// copyrights Fawad Haider
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 ;
  assign n6239 = x127 & x255 ;
  assign n6238 = x126 & x254 ;
  assign n6243 = n6239 ^ n6238 ;
  assign n6232 = x125 & x253 ;
  assign n6231 = x124 & x252 ;
  assign n6236 = n6232 ^ n6231 ;
  assign n6257 = n6243 ^ n6236 ;
  assign n6207 = x123 & x251 ;
  assign n6206 = x122 & x250 ;
  assign n6211 = n6207 ^ n6206 ;
  assign n6200 = x121 & x249 ;
  assign n6199 = x120 & x248 ;
  assign n6204 = n6200 ^ n6199 ;
  assign n6225 = n6211 ^ n6204 ;
  assign n6306 = n6257 ^ n6225 ;
  assign n6120 = x119 & x247 ;
  assign n6119 = x118 & x246 ;
  assign n6124 = n6120 ^ n6119 ;
  assign n6113 = x117 & x245 ;
  assign n6112 = x116 & x244 ;
  assign n6117 = n6113 ^ n6112 ;
  assign n6138 = n6124 ^ n6117 ;
  assign n6088 = x115 & x243 ;
  assign n6087 = x114 & x242 ;
  assign n6092 = n6088 ^ n6087 ;
  assign n6081 = x113 & x241 ;
  assign n6080 = x112 & x240 ;
  assign n6085 = n6081 ^ n6080 ;
  assign n6106 = n6092 ^ n6085 ;
  assign n6187 = n6138 ^ n6106 ;
  assign n6460 = n6306 ^ n6187 ;
  assign n5835 = x111 & x239 ;
  assign n5834 = x110 & x238 ;
  assign n5839 = n5835 ^ n5834 ;
  assign n5828 = x109 & x237 ;
  assign n5827 = x108 & x236 ;
  assign n5832 = n5828 ^ n5827 ;
  assign n5853 = n5839 ^ n5832 ;
  assign n5803 = x107 & x235 ;
  assign n5802 = x106 & x234 ;
  assign n5807 = n5803 ^ n5802 ;
  assign n5796 = x105 & x233 ;
  assign n5795 = x104 & x232 ;
  assign n5800 = n5796 ^ n5795 ;
  assign n5821 = n5807 ^ n5800 ;
  assign n5902 = n5853 ^ n5821 ;
  assign n5716 = x103 & x231 ;
  assign n5715 = x102 & x230 ;
  assign n5720 = n5716 ^ n5715 ;
  assign n5709 = x101 & x229 ;
  assign n5708 = x100 & x228 ;
  assign n5713 = n5709 ^ n5708 ;
  assign n5734 = n5720 ^ n5713 ;
  assign n5684 = x99 & x227 ;
  assign n5683 = x98 & x226 ;
  assign n5688 = n5684 ^ n5683 ;
  assign n5677 = x97 & x225 ;
  assign n5676 = x96 & x224 ;
  assign n5681 = n5677 ^ n5676 ;
  assign n5702 = n5688 ^ n5681 ;
  assign n5783 = n5734 ^ n5702 ;
  assign n6056 = n5902 ^ n5783 ;
  assign n6935 = n6460 ^ n6056 ;
  assign n4932 = x95 & x223 ;
  assign n4931 = x94 & x222 ;
  assign n4936 = n4932 ^ n4931 ;
  assign n4925 = x93 & x221 ;
  assign n4924 = x92 & x220 ;
  assign n4929 = n4925 ^ n4924 ;
  assign n4950 = n4936 ^ n4929 ;
  assign n4900 = x91 & x219 ;
  assign n4899 = x90 & x218 ;
  assign n4904 = n4900 ^ n4899 ;
  assign n4893 = x89 & x217 ;
  assign n4892 = x88 & x216 ;
  assign n4897 = n4893 ^ n4892 ;
  assign n4918 = n4904 ^ n4897 ;
  assign n4999 = n4950 ^ n4918 ;
  assign n4813 = x87 & x215 ;
  assign n4812 = x86 & x214 ;
  assign n4817 = n4813 ^ n4812 ;
  assign n4806 = x85 & x213 ;
  assign n4805 = x84 & x212 ;
  assign n4810 = n4806 ^ n4805 ;
  assign n4831 = n4817 ^ n4810 ;
  assign n4781 = x83 & x211 ;
  assign n4780 = x82 & x210 ;
  assign n4785 = n4781 ^ n4780 ;
  assign n4774 = x81 & x209 ;
  assign n4773 = x80 & x208 ;
  assign n4778 = n4774 ^ n4773 ;
  assign n4799 = n4785 ^ n4778 ;
  assign n4880 = n4831 ^ n4799 ;
  assign n5153 = n4999 ^ n4880 ;
  assign n4528 = x79 & x207 ;
  assign n4527 = x78 & x206 ;
  assign n4532 = n4528 ^ n4527 ;
  assign n4521 = x77 & x205 ;
  assign n4520 = x76 & x204 ;
  assign n4525 = n4521 ^ n4520 ;
  assign n4546 = n4532 ^ n4525 ;
  assign n4496 = x75 & x203 ;
  assign n4495 = x74 & x202 ;
  assign n4500 = n4496 ^ n4495 ;
  assign n4489 = x73 & x201 ;
  assign n4488 = x72 & x200 ;
  assign n4493 = n4489 ^ n4488 ;
  assign n4514 = n4500 ^ n4493 ;
  assign n4595 = n4546 ^ n4514 ;
  assign n4409 = x71 & x199 ;
  assign n4408 = x70 & x198 ;
  assign n4413 = n4409 ^ n4408 ;
  assign n4402 = x69 & x197 ;
  assign n4401 = x68 & x196 ;
  assign n4406 = n4402 ^ n4401 ;
  assign n4427 = n4413 ^ n4406 ;
  assign n4377 = x67 & x195 ;
  assign n4376 = x66 & x194 ;
  assign n4381 = n4377 ^ n4376 ;
  assign n4370 = x65 & x193 ;
  assign n4369 = x64 & x192 ;
  assign n4374 = n4370 ^ n4369 ;
  assign n4395 = n4381 ^ n4374 ;
  assign n4476 = n4427 ^ n4395 ;
  assign n4749 = n4595 ^ n4476 ;
  assign n5628 = n5153 ^ n4749 ;
  assign n8385 = n6935 ^ n5628 ;
  assign n2127 = x63 & x191 ;
  assign n2126 = x62 & x190 ;
  assign n2131 = n2127 ^ n2126 ;
  assign n2120 = x61 & x189 ;
  assign n2119 = x60 & x188 ;
  assign n2124 = n2120 ^ n2119 ;
  assign n2145 = n2131 ^ n2124 ;
  assign n2095 = x59 & x187 ;
  assign n2094 = x58 & x186 ;
  assign n2099 = n2095 ^ n2094 ;
  assign n2088 = x57 & x185 ;
  assign n2087 = x56 & x184 ;
  assign n2092 = n2088 ^ n2087 ;
  assign n2113 = n2099 ^ n2092 ;
  assign n2194 = n2145 ^ n2113 ;
  assign n2008 = x55 & x183 ;
  assign n2007 = x54 & x182 ;
  assign n2012 = n2008 ^ n2007 ;
  assign n2001 = x53 & x181 ;
  assign n2000 = x52 & x180 ;
  assign n2005 = n2001 ^ n2000 ;
  assign n2026 = n2012 ^ n2005 ;
  assign n1976 = x51 & x179 ;
  assign n1975 = x50 & x178 ;
  assign n1980 = n1976 ^ n1975 ;
  assign n1969 = x49 & x177 ;
  assign n1968 = x48 & x176 ;
  assign n1973 = n1969 ^ n1968 ;
  assign n1994 = n1980 ^ n1973 ;
  assign n2075 = n2026 ^ n1994 ;
  assign n2348 = n2194 ^ n2075 ;
  assign n1723 = x47 & x175 ;
  assign n1722 = x46 & x174 ;
  assign n1727 = n1723 ^ n1722 ;
  assign n1716 = x45 & x173 ;
  assign n1715 = x44 & x172 ;
  assign n1720 = n1716 ^ n1715 ;
  assign n1741 = n1727 ^ n1720 ;
  assign n1691 = x43 & x171 ;
  assign n1690 = x42 & x170 ;
  assign n1695 = n1691 ^ n1690 ;
  assign n1684 = x41 & x169 ;
  assign n1683 = x40 & x168 ;
  assign n1688 = n1684 ^ n1683 ;
  assign n1709 = n1695 ^ n1688 ;
  assign n1790 = n1741 ^ n1709 ;
  assign n1604 = x39 & x167 ;
  assign n1603 = x38 & x166 ;
  assign n1608 = n1604 ^ n1603 ;
  assign n1597 = x37 & x165 ;
  assign n1596 = x36 & x164 ;
  assign n1601 = n1597 ^ n1596 ;
  assign n1622 = n1608 ^ n1601 ;
  assign n1572 = x35 & x163 ;
  assign n1571 = x34 & x162 ;
  assign n1576 = n1572 ^ n1571 ;
  assign n1565 = x33 & x161 ;
  assign n1564 = x32 & x160 ;
  assign n1569 = n1565 ^ n1564 ;
  assign n1590 = n1576 ^ n1569 ;
  assign n1671 = n1622 ^ n1590 ;
  assign n1944 = n1790 ^ n1671 ;
  assign n2823 = n2348 ^ n1944 ;
  assign n820 = x31 & x159 ;
  assign n819 = x30 & x158 ;
  assign n824 = n820 ^ n819 ;
  assign n813 = x29 & x157 ;
  assign n812 = x28 & x156 ;
  assign n817 = n813 ^ n812 ;
  assign n838 = n824 ^ n817 ;
  assign n788 = x27 & x155 ;
  assign n787 = x26 & x154 ;
  assign n792 = n788 ^ n787 ;
  assign n781 = x25 & x153 ;
  assign n780 = x24 & x152 ;
  assign n785 = n781 ^ n780 ;
  assign n806 = n792 ^ n785 ;
  assign n887 = n838 ^ n806 ;
  assign n701 = x23 & x151 ;
  assign n700 = x22 & x150 ;
  assign n705 = n701 ^ n700 ;
  assign n694 = x21 & x149 ;
  assign n693 = x20 & x148 ;
  assign n698 = n694 ^ n693 ;
  assign n719 = n705 ^ n698 ;
  assign n669 = x19 & x147 ;
  assign n668 = x18 & x146 ;
  assign n673 = n669 ^ n668 ;
  assign n662 = x17 & x145 ;
  assign n661 = x16 & x144 ;
  assign n666 = n662 ^ n661 ;
  assign n687 = n673 ^ n666 ;
  assign n768 = n719 ^ n687 ;
  assign n1041 = n887 ^ n768 ;
  assign n416 = x15 & x143 ;
  assign n415 = x14 & x142 ;
  assign n420 = n416 ^ n415 ;
  assign n409 = x13 & x141 ;
  assign n408 = x12 & x140 ;
  assign n413 = n409 ^ n408 ;
  assign n434 = n420 ^ n413 ;
  assign n384 = x11 & x139 ;
  assign n383 = x10 & x138 ;
  assign n388 = n384 ^ n383 ;
  assign n377 = x9 & x137 ;
  assign n376 = x8 & x136 ;
  assign n381 = n377 ^ n376 ;
  assign n402 = n388 ^ n381 ;
  assign n483 = n434 ^ n402 ;
  assign n297 = x7 & x135 ;
  assign n296 = x6 & x134 ;
  assign n301 = n297 ^ n296 ;
  assign n290 = x5 & x133 ;
  assign n289 = x4 & x132 ;
  assign n294 = n290 ^ n289 ;
  assign n315 = n301 ^ n294 ;
  assign n265 = x3 & x131 ;
  assign n264 = x2 & x130 ;
  assign n269 = n265 ^ n264 ;
  assign n258 = x1 & x129 ;
  assign n257 = x0 & x128 ;
  assign n262 = n258 ^ n257 ;
  assign n283 = n269 ^ n262 ;
  assign n364 = n315 ^ n283 ;
  assign n637 = n483 ^ n364 ;
  assign n1516 = n1041 ^ n637 ;
  assign n4273 = n2823 ^ n1516 ;
  assign n12784 = n8385 ^ n4273 ;
  assign n6240 = x127 ^ x126 ;
  assign n6241 = x255 ^ x254 ;
  assign n6242 = n6240 & n6241 ;
  assign n6244 = n6242 ^ n6238 ;
  assign n6233 = x125 ^ x124 ;
  assign n6234 = x253 ^ x252 ;
  assign n6235 = n6233 & n6234 ;
  assign n6237 = n6235 ^ n6231 ;
  assign n6258 = n6244 ^ n6237 ;
  assign n6208 = x123 ^ x122 ;
  assign n6209 = x251 ^ x250 ;
  assign n6210 = n6208 & n6209 ;
  assign n6212 = n6210 ^ n6206 ;
  assign n6201 = x121 ^ x120 ;
  assign n6202 = x249 ^ x248 ;
  assign n6203 = n6201 & n6202 ;
  assign n6205 = n6203 ^ n6199 ;
  assign n6226 = n6212 ^ n6205 ;
  assign n6307 = n6258 ^ n6226 ;
  assign n6121 = x119 ^ x118 ;
  assign n6122 = x247 ^ x246 ;
  assign n6123 = n6121 & n6122 ;
  assign n6125 = n6123 ^ n6119 ;
  assign n6114 = x117 ^ x116 ;
  assign n6115 = x245 ^ x244 ;
  assign n6116 = n6114 & n6115 ;
  assign n6118 = n6116 ^ n6112 ;
  assign n6139 = n6125 ^ n6118 ;
  assign n6089 = x115 ^ x114 ;
  assign n6090 = x243 ^ x242 ;
  assign n6091 = n6089 & n6090 ;
  assign n6093 = n6091 ^ n6087 ;
  assign n6082 = x113 ^ x112 ;
  assign n6083 = x241 ^ x240 ;
  assign n6084 = n6082 & n6083 ;
  assign n6086 = n6084 ^ n6080 ;
  assign n6107 = n6093 ^ n6086 ;
  assign n6188 = n6139 ^ n6107 ;
  assign n6461 = n6307 ^ n6188 ;
  assign n5836 = x111 ^ x110 ;
  assign n5837 = x239 ^ x238 ;
  assign n5838 = n5836 & n5837 ;
  assign n5840 = n5838 ^ n5834 ;
  assign n5829 = x109 ^ x108 ;
  assign n5830 = x237 ^ x236 ;
  assign n5831 = n5829 & n5830 ;
  assign n5833 = n5831 ^ n5827 ;
  assign n5854 = n5840 ^ n5833 ;
  assign n5804 = x107 ^ x106 ;
  assign n5805 = x235 ^ x234 ;
  assign n5806 = n5804 & n5805 ;
  assign n5808 = n5806 ^ n5802 ;
  assign n5797 = x105 ^ x104 ;
  assign n5798 = x233 ^ x232 ;
  assign n5799 = n5797 & n5798 ;
  assign n5801 = n5799 ^ n5795 ;
  assign n5822 = n5808 ^ n5801 ;
  assign n5903 = n5854 ^ n5822 ;
  assign n5717 = x103 ^ x102 ;
  assign n5718 = x231 ^ x230 ;
  assign n5719 = n5717 & n5718 ;
  assign n5721 = n5719 ^ n5715 ;
  assign n5710 = x101 ^ x100 ;
  assign n5711 = x229 ^ x228 ;
  assign n5712 = n5710 & n5711 ;
  assign n5714 = n5712 ^ n5708 ;
  assign n5735 = n5721 ^ n5714 ;
  assign n5685 = x99 ^ x98 ;
  assign n5686 = x227 ^ x226 ;
  assign n5687 = n5685 & n5686 ;
  assign n5689 = n5687 ^ n5683 ;
  assign n5678 = x97 ^ x96 ;
  assign n5679 = x225 ^ x224 ;
  assign n5680 = n5678 & n5679 ;
  assign n5682 = n5680 ^ n5676 ;
  assign n5703 = n5689 ^ n5682 ;
  assign n5784 = n5735 ^ n5703 ;
  assign n6057 = n5903 ^ n5784 ;
  assign n6936 = n6461 ^ n6057 ;
  assign n4933 = x95 ^ x94 ;
  assign n4934 = x223 ^ x222 ;
  assign n4935 = n4933 & n4934 ;
  assign n4937 = n4935 ^ n4931 ;
  assign n4926 = x93 ^ x92 ;
  assign n4927 = x221 ^ x220 ;
  assign n4928 = n4926 & n4927 ;
  assign n4930 = n4928 ^ n4924 ;
  assign n4951 = n4937 ^ n4930 ;
  assign n4901 = x91 ^ x90 ;
  assign n4902 = x219 ^ x218 ;
  assign n4903 = n4901 & n4902 ;
  assign n4905 = n4903 ^ n4899 ;
  assign n4894 = x89 ^ x88 ;
  assign n4895 = x217 ^ x216 ;
  assign n4896 = n4894 & n4895 ;
  assign n4898 = n4896 ^ n4892 ;
  assign n4919 = n4905 ^ n4898 ;
  assign n5000 = n4951 ^ n4919 ;
  assign n4814 = x87 ^ x86 ;
  assign n4815 = x215 ^ x214 ;
  assign n4816 = n4814 & n4815 ;
  assign n4818 = n4816 ^ n4812 ;
  assign n4807 = x85 ^ x84 ;
  assign n4808 = x213 ^ x212 ;
  assign n4809 = n4807 & n4808 ;
  assign n4811 = n4809 ^ n4805 ;
  assign n4832 = n4818 ^ n4811 ;
  assign n4782 = x83 ^ x82 ;
  assign n4783 = x211 ^ x210 ;
  assign n4784 = n4782 & n4783 ;
  assign n4786 = n4784 ^ n4780 ;
  assign n4775 = x81 ^ x80 ;
  assign n4776 = x209 ^ x208 ;
  assign n4777 = n4775 & n4776 ;
  assign n4779 = n4777 ^ n4773 ;
  assign n4800 = n4786 ^ n4779 ;
  assign n4881 = n4832 ^ n4800 ;
  assign n5154 = n5000 ^ n4881 ;
  assign n4529 = x79 ^ x78 ;
  assign n4530 = x207 ^ x206 ;
  assign n4531 = n4529 & n4530 ;
  assign n4533 = n4531 ^ n4527 ;
  assign n4522 = x77 ^ x76 ;
  assign n4523 = x205 ^ x204 ;
  assign n4524 = n4522 & n4523 ;
  assign n4526 = n4524 ^ n4520 ;
  assign n4547 = n4533 ^ n4526 ;
  assign n4497 = x75 ^ x74 ;
  assign n4498 = x203 ^ x202 ;
  assign n4499 = n4497 & n4498 ;
  assign n4501 = n4499 ^ n4495 ;
  assign n4490 = x73 ^ x72 ;
  assign n4491 = x201 ^ x200 ;
  assign n4492 = n4490 & n4491 ;
  assign n4494 = n4492 ^ n4488 ;
  assign n4515 = n4501 ^ n4494 ;
  assign n4596 = n4547 ^ n4515 ;
  assign n4410 = x71 ^ x70 ;
  assign n4411 = x199 ^ x198 ;
  assign n4412 = n4410 & n4411 ;
  assign n4414 = n4412 ^ n4408 ;
  assign n4403 = x69 ^ x68 ;
  assign n4404 = x197 ^ x196 ;
  assign n4405 = n4403 & n4404 ;
  assign n4407 = n4405 ^ n4401 ;
  assign n4428 = n4414 ^ n4407 ;
  assign n4378 = x67 ^ x66 ;
  assign n4379 = x195 ^ x194 ;
  assign n4380 = n4378 & n4379 ;
  assign n4382 = n4380 ^ n4376 ;
  assign n4371 = x65 ^ x64 ;
  assign n4372 = x193 ^ x192 ;
  assign n4373 = n4371 & n4372 ;
  assign n4375 = n4373 ^ n4369 ;
  assign n4396 = n4382 ^ n4375 ;
  assign n4477 = n4428 ^ n4396 ;
  assign n4750 = n4596 ^ n4477 ;
  assign n5629 = n5154 ^ n4750 ;
  assign n8386 = n6936 ^ n5629 ;
  assign n2128 = x63 ^ x62 ;
  assign n2129 = x191 ^ x190 ;
  assign n2130 = n2128 & n2129 ;
  assign n2132 = n2130 ^ n2126 ;
  assign n2121 = x61 ^ x60 ;
  assign n2122 = x189 ^ x188 ;
  assign n2123 = n2121 & n2122 ;
  assign n2125 = n2123 ^ n2119 ;
  assign n2146 = n2132 ^ n2125 ;
  assign n2096 = x59 ^ x58 ;
  assign n2097 = x187 ^ x186 ;
  assign n2098 = n2096 & n2097 ;
  assign n2100 = n2098 ^ n2094 ;
  assign n2089 = x57 ^ x56 ;
  assign n2090 = x185 ^ x184 ;
  assign n2091 = n2089 & n2090 ;
  assign n2093 = n2091 ^ n2087 ;
  assign n2114 = n2100 ^ n2093 ;
  assign n2195 = n2146 ^ n2114 ;
  assign n2009 = x55 ^ x54 ;
  assign n2010 = x183 ^ x182 ;
  assign n2011 = n2009 & n2010 ;
  assign n2013 = n2011 ^ n2007 ;
  assign n2002 = x53 ^ x52 ;
  assign n2003 = x181 ^ x180 ;
  assign n2004 = n2002 & n2003 ;
  assign n2006 = n2004 ^ n2000 ;
  assign n2027 = n2013 ^ n2006 ;
  assign n1977 = x51 ^ x50 ;
  assign n1978 = x179 ^ x178 ;
  assign n1979 = n1977 & n1978 ;
  assign n1981 = n1979 ^ n1975 ;
  assign n1970 = x49 ^ x48 ;
  assign n1971 = x177 ^ x176 ;
  assign n1972 = n1970 & n1971 ;
  assign n1974 = n1972 ^ n1968 ;
  assign n1995 = n1981 ^ n1974 ;
  assign n2076 = n2027 ^ n1995 ;
  assign n2349 = n2195 ^ n2076 ;
  assign n1724 = x47 ^ x46 ;
  assign n1725 = x175 ^ x174 ;
  assign n1726 = n1724 & n1725 ;
  assign n1728 = n1726 ^ n1722 ;
  assign n1717 = x45 ^ x44 ;
  assign n1718 = x173 ^ x172 ;
  assign n1719 = n1717 & n1718 ;
  assign n1721 = n1719 ^ n1715 ;
  assign n1742 = n1728 ^ n1721 ;
  assign n1692 = x43 ^ x42 ;
  assign n1693 = x171 ^ x170 ;
  assign n1694 = n1692 & n1693 ;
  assign n1696 = n1694 ^ n1690 ;
  assign n1685 = x41 ^ x40 ;
  assign n1686 = x169 ^ x168 ;
  assign n1687 = n1685 & n1686 ;
  assign n1689 = n1687 ^ n1683 ;
  assign n1710 = n1696 ^ n1689 ;
  assign n1791 = n1742 ^ n1710 ;
  assign n1605 = x39 ^ x38 ;
  assign n1606 = x167 ^ x166 ;
  assign n1607 = n1605 & n1606 ;
  assign n1609 = n1607 ^ n1603 ;
  assign n1598 = x37 ^ x36 ;
  assign n1599 = x165 ^ x164 ;
  assign n1600 = n1598 & n1599 ;
  assign n1602 = n1600 ^ n1596 ;
  assign n1623 = n1609 ^ n1602 ;
  assign n1573 = x35 ^ x34 ;
  assign n1574 = x163 ^ x162 ;
  assign n1575 = n1573 & n1574 ;
  assign n1577 = n1575 ^ n1571 ;
  assign n1566 = x33 ^ x32 ;
  assign n1567 = x161 ^ x160 ;
  assign n1568 = n1566 & n1567 ;
  assign n1570 = n1568 ^ n1564 ;
  assign n1591 = n1577 ^ n1570 ;
  assign n1672 = n1623 ^ n1591 ;
  assign n1945 = n1791 ^ n1672 ;
  assign n2824 = n2349 ^ n1945 ;
  assign n821 = x31 ^ x30 ;
  assign n822 = x159 ^ x158 ;
  assign n823 = n821 & n822 ;
  assign n825 = n823 ^ n819 ;
  assign n814 = x29 ^ x28 ;
  assign n815 = x157 ^ x156 ;
  assign n816 = n814 & n815 ;
  assign n818 = n816 ^ n812 ;
  assign n839 = n825 ^ n818 ;
  assign n789 = x27 ^ x26 ;
  assign n790 = x155 ^ x154 ;
  assign n791 = n789 & n790 ;
  assign n793 = n791 ^ n787 ;
  assign n782 = x25 ^ x24 ;
  assign n783 = x153 ^ x152 ;
  assign n784 = n782 & n783 ;
  assign n786 = n784 ^ n780 ;
  assign n807 = n793 ^ n786 ;
  assign n888 = n839 ^ n807 ;
  assign n702 = x23 ^ x22 ;
  assign n703 = x151 ^ x150 ;
  assign n704 = n702 & n703 ;
  assign n706 = n704 ^ n700 ;
  assign n695 = x21 ^ x20 ;
  assign n696 = x149 ^ x148 ;
  assign n697 = n695 & n696 ;
  assign n699 = n697 ^ n693 ;
  assign n720 = n706 ^ n699 ;
  assign n670 = x19 ^ x18 ;
  assign n671 = x147 ^ x146 ;
  assign n672 = n670 & n671 ;
  assign n674 = n672 ^ n668 ;
  assign n663 = x17 ^ x16 ;
  assign n664 = x145 ^ x144 ;
  assign n665 = n663 & n664 ;
  assign n667 = n665 ^ n661 ;
  assign n688 = n674 ^ n667 ;
  assign n769 = n720 ^ n688 ;
  assign n1042 = n888 ^ n769 ;
  assign n417 = x15 ^ x14 ;
  assign n418 = x143 ^ x142 ;
  assign n419 = n417 & n418 ;
  assign n421 = n419 ^ n415 ;
  assign n410 = x13 ^ x12 ;
  assign n411 = x141 ^ x140 ;
  assign n412 = n410 & n411 ;
  assign n414 = n412 ^ n408 ;
  assign n435 = n421 ^ n414 ;
  assign n385 = x11 ^ x10 ;
  assign n386 = x139 ^ x138 ;
  assign n387 = n385 & n386 ;
  assign n389 = n387 ^ n383 ;
  assign n378 = x9 ^ x8 ;
  assign n379 = x137 ^ x136 ;
  assign n380 = n378 & n379 ;
  assign n382 = n380 ^ n376 ;
  assign n403 = n389 ^ n382 ;
  assign n484 = n435 ^ n403 ;
  assign n298 = x7 ^ x6 ;
  assign n299 = x135 ^ x134 ;
  assign n300 = n298 & n299 ;
  assign n302 = n300 ^ n296 ;
  assign n291 = x5 ^ x4 ;
  assign n292 = x133 ^ x132 ;
  assign n293 = n291 & n292 ;
  assign n295 = n293 ^ n289 ;
  assign n316 = n302 ^ n295 ;
  assign n266 = x3 ^ x2 ;
  assign n267 = x131 ^ x130 ;
  assign n268 = n266 & n267 ;
  assign n270 = n268 ^ n264 ;
  assign n259 = x1 ^ x0 ;
  assign n260 = x129 ^ x128 ;
  assign n261 = n259 & n260 ;
  assign n263 = n261 ^ n257 ;
  assign n284 = n270 ^ n263 ;
  assign n365 = n316 ^ n284 ;
  assign n638 = n484 ^ n365 ;
  assign n1517 = n1042 ^ n638 ;
  assign n4274 = n2824 ^ n1517 ;
  assign n12785 = n8386 ^ n4274 ;
  assign n6247 = x127 ^ x125 ;
  assign n6248 = x255 ^ x253 ;
  assign n6251 = n6247 & n6248 ;
  assign n6245 = x126 ^ x124 ;
  assign n6246 = x254 ^ x252 ;
  assign n6250 = n6245 & n6246 ;
  assign n6255 = n6251 ^ n6250 ;
  assign n6259 = n6257 ^ n6255 ;
  assign n6260 = n6259 ^ n6244 ;
  assign n6215 = x123 ^ x121 ;
  assign n6216 = x251 ^ x249 ;
  assign n6219 = n6215 & n6216 ;
  assign n6213 = x122 ^ x120 ;
  assign n6214 = x250 ^ x248 ;
  assign n6218 = n6213 & n6214 ;
  assign n6223 = n6219 ^ n6218 ;
  assign n6227 = n6225 ^ n6223 ;
  assign n6228 = n6227 ^ n6212 ;
  assign n6308 = n6260 ^ n6228 ;
  assign n6128 = x119 ^ x117 ;
  assign n6129 = x247 ^ x245 ;
  assign n6132 = n6128 & n6129 ;
  assign n6126 = x118 ^ x116 ;
  assign n6127 = x246 ^ x244 ;
  assign n6131 = n6126 & n6127 ;
  assign n6136 = n6132 ^ n6131 ;
  assign n6140 = n6138 ^ n6136 ;
  assign n6141 = n6140 ^ n6125 ;
  assign n6096 = x115 ^ x113 ;
  assign n6097 = x243 ^ x241 ;
  assign n6100 = n6096 & n6097 ;
  assign n6094 = x114 ^ x112 ;
  assign n6095 = x242 ^ x240 ;
  assign n6099 = n6094 & n6095 ;
  assign n6104 = n6100 ^ n6099 ;
  assign n6108 = n6106 ^ n6104 ;
  assign n6109 = n6108 ^ n6093 ;
  assign n6189 = n6141 ^ n6109 ;
  assign n6462 = n6308 ^ n6189 ;
  assign n5843 = x111 ^ x109 ;
  assign n5844 = x239 ^ x237 ;
  assign n5847 = n5843 & n5844 ;
  assign n5841 = x110 ^ x108 ;
  assign n5842 = x238 ^ x236 ;
  assign n5846 = n5841 & n5842 ;
  assign n5851 = n5847 ^ n5846 ;
  assign n5855 = n5853 ^ n5851 ;
  assign n5856 = n5855 ^ n5840 ;
  assign n5811 = x107 ^ x105 ;
  assign n5812 = x235 ^ x233 ;
  assign n5815 = n5811 & n5812 ;
  assign n5809 = x106 ^ x104 ;
  assign n5810 = x234 ^ x232 ;
  assign n5814 = n5809 & n5810 ;
  assign n5819 = n5815 ^ n5814 ;
  assign n5823 = n5821 ^ n5819 ;
  assign n5824 = n5823 ^ n5808 ;
  assign n5904 = n5856 ^ n5824 ;
  assign n5724 = x103 ^ x101 ;
  assign n5725 = x231 ^ x229 ;
  assign n5728 = n5724 & n5725 ;
  assign n5722 = x102 ^ x100 ;
  assign n5723 = x230 ^ x228 ;
  assign n5727 = n5722 & n5723 ;
  assign n5732 = n5728 ^ n5727 ;
  assign n5736 = n5734 ^ n5732 ;
  assign n5737 = n5736 ^ n5721 ;
  assign n5692 = x99 ^ x97 ;
  assign n5693 = x227 ^ x225 ;
  assign n5696 = n5692 & n5693 ;
  assign n5690 = x98 ^ x96 ;
  assign n5691 = x226 ^ x224 ;
  assign n5695 = n5690 & n5691 ;
  assign n5700 = n5696 ^ n5695 ;
  assign n5704 = n5702 ^ n5700 ;
  assign n5705 = n5704 ^ n5689 ;
  assign n5785 = n5737 ^ n5705 ;
  assign n6058 = n5904 ^ n5785 ;
  assign n6937 = n6462 ^ n6058 ;
  assign n4940 = x95 ^ x93 ;
  assign n4941 = x223 ^ x221 ;
  assign n4944 = n4940 & n4941 ;
  assign n4938 = x94 ^ x92 ;
  assign n4939 = x222 ^ x220 ;
  assign n4943 = n4938 & n4939 ;
  assign n4948 = n4944 ^ n4943 ;
  assign n4952 = n4950 ^ n4948 ;
  assign n4953 = n4952 ^ n4937 ;
  assign n4908 = x91 ^ x89 ;
  assign n4909 = x219 ^ x217 ;
  assign n4912 = n4908 & n4909 ;
  assign n4906 = x90 ^ x88 ;
  assign n4907 = x218 ^ x216 ;
  assign n4911 = n4906 & n4907 ;
  assign n4916 = n4912 ^ n4911 ;
  assign n4920 = n4918 ^ n4916 ;
  assign n4921 = n4920 ^ n4905 ;
  assign n5001 = n4953 ^ n4921 ;
  assign n4821 = x87 ^ x85 ;
  assign n4822 = x215 ^ x213 ;
  assign n4825 = n4821 & n4822 ;
  assign n4819 = x86 ^ x84 ;
  assign n4820 = x214 ^ x212 ;
  assign n4824 = n4819 & n4820 ;
  assign n4829 = n4825 ^ n4824 ;
  assign n4833 = n4831 ^ n4829 ;
  assign n4834 = n4833 ^ n4818 ;
  assign n4789 = x83 ^ x81 ;
  assign n4790 = x211 ^ x209 ;
  assign n4793 = n4789 & n4790 ;
  assign n4787 = x82 ^ x80 ;
  assign n4788 = x210 ^ x208 ;
  assign n4792 = n4787 & n4788 ;
  assign n4797 = n4793 ^ n4792 ;
  assign n4801 = n4799 ^ n4797 ;
  assign n4802 = n4801 ^ n4786 ;
  assign n4882 = n4834 ^ n4802 ;
  assign n5155 = n5001 ^ n4882 ;
  assign n4536 = x79 ^ x77 ;
  assign n4537 = x207 ^ x205 ;
  assign n4540 = n4536 & n4537 ;
  assign n4534 = x78 ^ x76 ;
  assign n4535 = x206 ^ x204 ;
  assign n4539 = n4534 & n4535 ;
  assign n4544 = n4540 ^ n4539 ;
  assign n4548 = n4546 ^ n4544 ;
  assign n4549 = n4548 ^ n4533 ;
  assign n4504 = x75 ^ x73 ;
  assign n4505 = x203 ^ x201 ;
  assign n4508 = n4504 & n4505 ;
  assign n4502 = x74 ^ x72 ;
  assign n4503 = x202 ^ x200 ;
  assign n4507 = n4502 & n4503 ;
  assign n4512 = n4508 ^ n4507 ;
  assign n4516 = n4514 ^ n4512 ;
  assign n4517 = n4516 ^ n4501 ;
  assign n4597 = n4549 ^ n4517 ;
  assign n4417 = x71 ^ x69 ;
  assign n4418 = x199 ^ x197 ;
  assign n4421 = n4417 & n4418 ;
  assign n4415 = x70 ^ x68 ;
  assign n4416 = x198 ^ x196 ;
  assign n4420 = n4415 & n4416 ;
  assign n4425 = n4421 ^ n4420 ;
  assign n4429 = n4427 ^ n4425 ;
  assign n4430 = n4429 ^ n4414 ;
  assign n4385 = x67 ^ x65 ;
  assign n4386 = x195 ^ x193 ;
  assign n4389 = n4385 & n4386 ;
  assign n4383 = x66 ^ x64 ;
  assign n4384 = x194 ^ x192 ;
  assign n4388 = n4383 & n4384 ;
  assign n4393 = n4389 ^ n4388 ;
  assign n4397 = n4395 ^ n4393 ;
  assign n4398 = n4397 ^ n4382 ;
  assign n4478 = n4430 ^ n4398 ;
  assign n4751 = n4597 ^ n4478 ;
  assign n5630 = n5155 ^ n4751 ;
  assign n8387 = n6937 ^ n5630 ;
  assign n2135 = x63 ^ x61 ;
  assign n2136 = x191 ^ x189 ;
  assign n2139 = n2135 & n2136 ;
  assign n2133 = x62 ^ x60 ;
  assign n2134 = x190 ^ x188 ;
  assign n2138 = n2133 & n2134 ;
  assign n2143 = n2139 ^ n2138 ;
  assign n2147 = n2145 ^ n2143 ;
  assign n2148 = n2147 ^ n2132 ;
  assign n2103 = x59 ^ x57 ;
  assign n2104 = x187 ^ x185 ;
  assign n2107 = n2103 & n2104 ;
  assign n2101 = x58 ^ x56 ;
  assign n2102 = x186 ^ x184 ;
  assign n2106 = n2101 & n2102 ;
  assign n2111 = n2107 ^ n2106 ;
  assign n2115 = n2113 ^ n2111 ;
  assign n2116 = n2115 ^ n2100 ;
  assign n2196 = n2148 ^ n2116 ;
  assign n2016 = x55 ^ x53 ;
  assign n2017 = x183 ^ x181 ;
  assign n2020 = n2016 & n2017 ;
  assign n2014 = x54 ^ x52 ;
  assign n2015 = x182 ^ x180 ;
  assign n2019 = n2014 & n2015 ;
  assign n2024 = n2020 ^ n2019 ;
  assign n2028 = n2026 ^ n2024 ;
  assign n2029 = n2028 ^ n2013 ;
  assign n1984 = x51 ^ x49 ;
  assign n1985 = x179 ^ x177 ;
  assign n1988 = n1984 & n1985 ;
  assign n1982 = x50 ^ x48 ;
  assign n1983 = x178 ^ x176 ;
  assign n1987 = n1982 & n1983 ;
  assign n1992 = n1988 ^ n1987 ;
  assign n1996 = n1994 ^ n1992 ;
  assign n1997 = n1996 ^ n1981 ;
  assign n2077 = n2029 ^ n1997 ;
  assign n2350 = n2196 ^ n2077 ;
  assign n1731 = x47 ^ x45 ;
  assign n1732 = x175 ^ x173 ;
  assign n1735 = n1731 & n1732 ;
  assign n1729 = x46 ^ x44 ;
  assign n1730 = x174 ^ x172 ;
  assign n1734 = n1729 & n1730 ;
  assign n1739 = n1735 ^ n1734 ;
  assign n1743 = n1741 ^ n1739 ;
  assign n1744 = n1743 ^ n1728 ;
  assign n1699 = x43 ^ x41 ;
  assign n1700 = x171 ^ x169 ;
  assign n1703 = n1699 & n1700 ;
  assign n1697 = x42 ^ x40 ;
  assign n1698 = x170 ^ x168 ;
  assign n1702 = n1697 & n1698 ;
  assign n1707 = n1703 ^ n1702 ;
  assign n1711 = n1709 ^ n1707 ;
  assign n1712 = n1711 ^ n1696 ;
  assign n1792 = n1744 ^ n1712 ;
  assign n1612 = x39 ^ x37 ;
  assign n1613 = x167 ^ x165 ;
  assign n1616 = n1612 & n1613 ;
  assign n1610 = x38 ^ x36 ;
  assign n1611 = x166 ^ x164 ;
  assign n1615 = n1610 & n1611 ;
  assign n1620 = n1616 ^ n1615 ;
  assign n1624 = n1622 ^ n1620 ;
  assign n1625 = n1624 ^ n1609 ;
  assign n1580 = x35 ^ x33 ;
  assign n1581 = x163 ^ x161 ;
  assign n1584 = n1580 & n1581 ;
  assign n1578 = x34 ^ x32 ;
  assign n1579 = x162 ^ x160 ;
  assign n1583 = n1578 & n1579 ;
  assign n1588 = n1584 ^ n1583 ;
  assign n1592 = n1590 ^ n1588 ;
  assign n1593 = n1592 ^ n1577 ;
  assign n1673 = n1625 ^ n1593 ;
  assign n1946 = n1792 ^ n1673 ;
  assign n2825 = n2350 ^ n1946 ;
  assign n828 = x31 ^ x29 ;
  assign n829 = x159 ^ x157 ;
  assign n832 = n828 & n829 ;
  assign n826 = x30 ^ x28 ;
  assign n827 = x158 ^ x156 ;
  assign n831 = n826 & n827 ;
  assign n836 = n832 ^ n831 ;
  assign n840 = n838 ^ n836 ;
  assign n841 = n840 ^ n825 ;
  assign n796 = x27 ^ x25 ;
  assign n797 = x155 ^ x153 ;
  assign n800 = n796 & n797 ;
  assign n794 = x26 ^ x24 ;
  assign n795 = x154 ^ x152 ;
  assign n799 = n794 & n795 ;
  assign n804 = n800 ^ n799 ;
  assign n808 = n806 ^ n804 ;
  assign n809 = n808 ^ n793 ;
  assign n889 = n841 ^ n809 ;
  assign n709 = x23 ^ x21 ;
  assign n710 = x151 ^ x149 ;
  assign n713 = n709 & n710 ;
  assign n707 = x22 ^ x20 ;
  assign n708 = x150 ^ x148 ;
  assign n712 = n707 & n708 ;
  assign n717 = n713 ^ n712 ;
  assign n721 = n719 ^ n717 ;
  assign n722 = n721 ^ n706 ;
  assign n677 = x19 ^ x17 ;
  assign n678 = x147 ^ x145 ;
  assign n681 = n677 & n678 ;
  assign n675 = x18 ^ x16 ;
  assign n676 = x146 ^ x144 ;
  assign n680 = n675 & n676 ;
  assign n685 = n681 ^ n680 ;
  assign n689 = n687 ^ n685 ;
  assign n690 = n689 ^ n674 ;
  assign n770 = n722 ^ n690 ;
  assign n1043 = n889 ^ n770 ;
  assign n424 = x15 ^ x13 ;
  assign n425 = x143 ^ x141 ;
  assign n428 = n424 & n425 ;
  assign n422 = x14 ^ x12 ;
  assign n423 = x142 ^ x140 ;
  assign n427 = n422 & n423 ;
  assign n432 = n428 ^ n427 ;
  assign n436 = n434 ^ n432 ;
  assign n437 = n436 ^ n421 ;
  assign n392 = x11 ^ x9 ;
  assign n393 = x139 ^ x137 ;
  assign n396 = n392 & n393 ;
  assign n390 = x10 ^ x8 ;
  assign n391 = x138 ^ x136 ;
  assign n395 = n390 & n391 ;
  assign n400 = n396 ^ n395 ;
  assign n404 = n402 ^ n400 ;
  assign n405 = n404 ^ n389 ;
  assign n485 = n437 ^ n405 ;
  assign n305 = x7 ^ x5 ;
  assign n306 = x135 ^ x133 ;
  assign n309 = n305 & n306 ;
  assign n303 = x6 ^ x4 ;
  assign n304 = x134 ^ x132 ;
  assign n308 = n303 & n304 ;
  assign n313 = n309 ^ n308 ;
  assign n317 = n315 ^ n313 ;
  assign n318 = n317 ^ n302 ;
  assign n273 = x3 ^ x1 ;
  assign n274 = x131 ^ x129 ;
  assign n277 = n273 & n274 ;
  assign n271 = x2 ^ x0 ;
  assign n272 = x130 ^ x128 ;
  assign n276 = n271 & n272 ;
  assign n281 = n277 ^ n276 ;
  assign n285 = n283 ^ n281 ;
  assign n286 = n285 ^ n270 ;
  assign n366 = n318 ^ n286 ;
  assign n639 = n485 ^ n366 ;
  assign n1518 = n1043 ^ n639 ;
  assign n4275 = n2825 ^ n1518 ;
  assign n12786 = n8387 ^ n4275 ;
  assign n6252 = n6247 ^ n6245 ;
  assign n6253 = n6248 ^ n6246 ;
  assign n6254 = n6252 & n6253 ;
  assign n6256 = n6254 ^ n6250 ;
  assign n6261 = n6258 ^ n6256 ;
  assign n6249 = n6244 ^ n6243 ;
  assign n6262 = n6261 ^ n6249 ;
  assign n6220 = n6215 ^ n6213 ;
  assign n6221 = n6216 ^ n6214 ;
  assign n6222 = n6220 & n6221 ;
  assign n6224 = n6222 ^ n6218 ;
  assign n6229 = n6226 ^ n6224 ;
  assign n6217 = n6212 ^ n6211 ;
  assign n6230 = n6229 ^ n6217 ;
  assign n6309 = n6262 ^ n6230 ;
  assign n6133 = n6128 ^ n6126 ;
  assign n6134 = n6129 ^ n6127 ;
  assign n6135 = n6133 & n6134 ;
  assign n6137 = n6135 ^ n6131 ;
  assign n6142 = n6139 ^ n6137 ;
  assign n6130 = n6125 ^ n6124 ;
  assign n6143 = n6142 ^ n6130 ;
  assign n6101 = n6096 ^ n6094 ;
  assign n6102 = n6097 ^ n6095 ;
  assign n6103 = n6101 & n6102 ;
  assign n6105 = n6103 ^ n6099 ;
  assign n6110 = n6107 ^ n6105 ;
  assign n6098 = n6093 ^ n6092 ;
  assign n6111 = n6110 ^ n6098 ;
  assign n6190 = n6143 ^ n6111 ;
  assign n6463 = n6309 ^ n6190 ;
  assign n5848 = n5843 ^ n5841 ;
  assign n5849 = n5844 ^ n5842 ;
  assign n5850 = n5848 & n5849 ;
  assign n5852 = n5850 ^ n5846 ;
  assign n5857 = n5854 ^ n5852 ;
  assign n5845 = n5840 ^ n5839 ;
  assign n5858 = n5857 ^ n5845 ;
  assign n5816 = n5811 ^ n5809 ;
  assign n5817 = n5812 ^ n5810 ;
  assign n5818 = n5816 & n5817 ;
  assign n5820 = n5818 ^ n5814 ;
  assign n5825 = n5822 ^ n5820 ;
  assign n5813 = n5808 ^ n5807 ;
  assign n5826 = n5825 ^ n5813 ;
  assign n5905 = n5858 ^ n5826 ;
  assign n5729 = n5724 ^ n5722 ;
  assign n5730 = n5725 ^ n5723 ;
  assign n5731 = n5729 & n5730 ;
  assign n5733 = n5731 ^ n5727 ;
  assign n5738 = n5735 ^ n5733 ;
  assign n5726 = n5721 ^ n5720 ;
  assign n5739 = n5738 ^ n5726 ;
  assign n5697 = n5692 ^ n5690 ;
  assign n5698 = n5693 ^ n5691 ;
  assign n5699 = n5697 & n5698 ;
  assign n5701 = n5699 ^ n5695 ;
  assign n5706 = n5703 ^ n5701 ;
  assign n5694 = n5689 ^ n5688 ;
  assign n5707 = n5706 ^ n5694 ;
  assign n5786 = n5739 ^ n5707 ;
  assign n6059 = n5905 ^ n5786 ;
  assign n6938 = n6463 ^ n6059 ;
  assign n4945 = n4940 ^ n4938 ;
  assign n4946 = n4941 ^ n4939 ;
  assign n4947 = n4945 & n4946 ;
  assign n4949 = n4947 ^ n4943 ;
  assign n4954 = n4951 ^ n4949 ;
  assign n4942 = n4937 ^ n4936 ;
  assign n4955 = n4954 ^ n4942 ;
  assign n4913 = n4908 ^ n4906 ;
  assign n4914 = n4909 ^ n4907 ;
  assign n4915 = n4913 & n4914 ;
  assign n4917 = n4915 ^ n4911 ;
  assign n4922 = n4919 ^ n4917 ;
  assign n4910 = n4905 ^ n4904 ;
  assign n4923 = n4922 ^ n4910 ;
  assign n5002 = n4955 ^ n4923 ;
  assign n4826 = n4821 ^ n4819 ;
  assign n4827 = n4822 ^ n4820 ;
  assign n4828 = n4826 & n4827 ;
  assign n4830 = n4828 ^ n4824 ;
  assign n4835 = n4832 ^ n4830 ;
  assign n4823 = n4818 ^ n4817 ;
  assign n4836 = n4835 ^ n4823 ;
  assign n4794 = n4789 ^ n4787 ;
  assign n4795 = n4790 ^ n4788 ;
  assign n4796 = n4794 & n4795 ;
  assign n4798 = n4796 ^ n4792 ;
  assign n4803 = n4800 ^ n4798 ;
  assign n4791 = n4786 ^ n4785 ;
  assign n4804 = n4803 ^ n4791 ;
  assign n4883 = n4836 ^ n4804 ;
  assign n5156 = n5002 ^ n4883 ;
  assign n4541 = n4536 ^ n4534 ;
  assign n4542 = n4537 ^ n4535 ;
  assign n4543 = n4541 & n4542 ;
  assign n4545 = n4543 ^ n4539 ;
  assign n4550 = n4547 ^ n4545 ;
  assign n4538 = n4533 ^ n4532 ;
  assign n4551 = n4550 ^ n4538 ;
  assign n4509 = n4504 ^ n4502 ;
  assign n4510 = n4505 ^ n4503 ;
  assign n4511 = n4509 & n4510 ;
  assign n4513 = n4511 ^ n4507 ;
  assign n4518 = n4515 ^ n4513 ;
  assign n4506 = n4501 ^ n4500 ;
  assign n4519 = n4518 ^ n4506 ;
  assign n4598 = n4551 ^ n4519 ;
  assign n4422 = n4417 ^ n4415 ;
  assign n4423 = n4418 ^ n4416 ;
  assign n4424 = n4422 & n4423 ;
  assign n4426 = n4424 ^ n4420 ;
  assign n4431 = n4428 ^ n4426 ;
  assign n4419 = n4414 ^ n4413 ;
  assign n4432 = n4431 ^ n4419 ;
  assign n4390 = n4385 ^ n4383 ;
  assign n4391 = n4386 ^ n4384 ;
  assign n4392 = n4390 & n4391 ;
  assign n4394 = n4392 ^ n4388 ;
  assign n4399 = n4396 ^ n4394 ;
  assign n4387 = n4382 ^ n4381 ;
  assign n4400 = n4399 ^ n4387 ;
  assign n4479 = n4432 ^ n4400 ;
  assign n4752 = n4598 ^ n4479 ;
  assign n5631 = n5156 ^ n4752 ;
  assign n8388 = n6938 ^ n5631 ;
  assign n2140 = n2135 ^ n2133 ;
  assign n2141 = n2136 ^ n2134 ;
  assign n2142 = n2140 & n2141 ;
  assign n2144 = n2142 ^ n2138 ;
  assign n2149 = n2146 ^ n2144 ;
  assign n2137 = n2132 ^ n2131 ;
  assign n2150 = n2149 ^ n2137 ;
  assign n2108 = n2103 ^ n2101 ;
  assign n2109 = n2104 ^ n2102 ;
  assign n2110 = n2108 & n2109 ;
  assign n2112 = n2110 ^ n2106 ;
  assign n2117 = n2114 ^ n2112 ;
  assign n2105 = n2100 ^ n2099 ;
  assign n2118 = n2117 ^ n2105 ;
  assign n2197 = n2150 ^ n2118 ;
  assign n2021 = n2016 ^ n2014 ;
  assign n2022 = n2017 ^ n2015 ;
  assign n2023 = n2021 & n2022 ;
  assign n2025 = n2023 ^ n2019 ;
  assign n2030 = n2027 ^ n2025 ;
  assign n2018 = n2013 ^ n2012 ;
  assign n2031 = n2030 ^ n2018 ;
  assign n1989 = n1984 ^ n1982 ;
  assign n1990 = n1985 ^ n1983 ;
  assign n1991 = n1989 & n1990 ;
  assign n1993 = n1991 ^ n1987 ;
  assign n1998 = n1995 ^ n1993 ;
  assign n1986 = n1981 ^ n1980 ;
  assign n1999 = n1998 ^ n1986 ;
  assign n2078 = n2031 ^ n1999 ;
  assign n2351 = n2197 ^ n2078 ;
  assign n1736 = n1731 ^ n1729 ;
  assign n1737 = n1732 ^ n1730 ;
  assign n1738 = n1736 & n1737 ;
  assign n1740 = n1738 ^ n1734 ;
  assign n1745 = n1742 ^ n1740 ;
  assign n1733 = n1728 ^ n1727 ;
  assign n1746 = n1745 ^ n1733 ;
  assign n1704 = n1699 ^ n1697 ;
  assign n1705 = n1700 ^ n1698 ;
  assign n1706 = n1704 & n1705 ;
  assign n1708 = n1706 ^ n1702 ;
  assign n1713 = n1710 ^ n1708 ;
  assign n1701 = n1696 ^ n1695 ;
  assign n1714 = n1713 ^ n1701 ;
  assign n1793 = n1746 ^ n1714 ;
  assign n1617 = n1612 ^ n1610 ;
  assign n1618 = n1613 ^ n1611 ;
  assign n1619 = n1617 & n1618 ;
  assign n1621 = n1619 ^ n1615 ;
  assign n1626 = n1623 ^ n1621 ;
  assign n1614 = n1609 ^ n1608 ;
  assign n1627 = n1626 ^ n1614 ;
  assign n1585 = n1580 ^ n1578 ;
  assign n1586 = n1581 ^ n1579 ;
  assign n1587 = n1585 & n1586 ;
  assign n1589 = n1587 ^ n1583 ;
  assign n1594 = n1591 ^ n1589 ;
  assign n1582 = n1577 ^ n1576 ;
  assign n1595 = n1594 ^ n1582 ;
  assign n1674 = n1627 ^ n1595 ;
  assign n1947 = n1793 ^ n1674 ;
  assign n2826 = n2351 ^ n1947 ;
  assign n833 = n828 ^ n826 ;
  assign n834 = n829 ^ n827 ;
  assign n835 = n833 & n834 ;
  assign n837 = n835 ^ n831 ;
  assign n842 = n839 ^ n837 ;
  assign n830 = n825 ^ n824 ;
  assign n843 = n842 ^ n830 ;
  assign n801 = n796 ^ n794 ;
  assign n802 = n797 ^ n795 ;
  assign n803 = n801 & n802 ;
  assign n805 = n803 ^ n799 ;
  assign n810 = n807 ^ n805 ;
  assign n798 = n793 ^ n792 ;
  assign n811 = n810 ^ n798 ;
  assign n890 = n843 ^ n811 ;
  assign n714 = n709 ^ n707 ;
  assign n715 = n710 ^ n708 ;
  assign n716 = n714 & n715 ;
  assign n718 = n716 ^ n712 ;
  assign n723 = n720 ^ n718 ;
  assign n711 = n706 ^ n705 ;
  assign n724 = n723 ^ n711 ;
  assign n682 = n677 ^ n675 ;
  assign n683 = n678 ^ n676 ;
  assign n684 = n682 & n683 ;
  assign n686 = n684 ^ n680 ;
  assign n691 = n688 ^ n686 ;
  assign n679 = n674 ^ n673 ;
  assign n692 = n691 ^ n679 ;
  assign n771 = n724 ^ n692 ;
  assign n1044 = n890 ^ n771 ;
  assign n429 = n424 ^ n422 ;
  assign n430 = n425 ^ n423 ;
  assign n431 = n429 & n430 ;
  assign n433 = n431 ^ n427 ;
  assign n438 = n435 ^ n433 ;
  assign n426 = n421 ^ n420 ;
  assign n439 = n438 ^ n426 ;
  assign n397 = n392 ^ n390 ;
  assign n398 = n393 ^ n391 ;
  assign n399 = n397 & n398 ;
  assign n401 = n399 ^ n395 ;
  assign n406 = n403 ^ n401 ;
  assign n394 = n389 ^ n388 ;
  assign n407 = n406 ^ n394 ;
  assign n486 = n439 ^ n407 ;
  assign n310 = n305 ^ n303 ;
  assign n311 = n306 ^ n304 ;
  assign n312 = n310 & n311 ;
  assign n314 = n312 ^ n308 ;
  assign n319 = n316 ^ n314 ;
  assign n307 = n302 ^ n301 ;
  assign n320 = n319 ^ n307 ;
  assign n278 = n273 ^ n271 ;
  assign n279 = n274 ^ n272 ;
  assign n280 = n278 & n279 ;
  assign n282 = n280 ^ n276 ;
  assign n287 = n284 ^ n282 ;
  assign n275 = n270 ^ n269 ;
  assign n288 = n287 ^ n275 ;
  assign n367 = n320 ^ n288 ;
  assign n640 = n486 ^ n367 ;
  assign n1519 = n1044 ^ n640 ;
  assign n4276 = n2826 ^ n1519 ;
  assign n12787 = n8388 ^ n4276 ;
  assign n6269 = x127 ^ x123 ;
  assign n6270 = x255 ^ x251 ;
  assign n6282 = n6269 & n6270 ;
  assign n6267 = x126 ^ x122 ;
  assign n6268 = x254 ^ x250 ;
  assign n6281 = n6267 & n6268 ;
  assign n6286 = n6282 ^ n6281 ;
  assign n6265 = x125 ^ x121 ;
  assign n6266 = x253 ^ x249 ;
  assign n6275 = n6265 & n6266 ;
  assign n6263 = x124 ^ x120 ;
  assign n6264 = x252 ^ x248 ;
  assign n6274 = n6263 & n6264 ;
  assign n6279 = n6275 ^ n6274 ;
  assign n6300 = n6286 ^ n6279 ;
  assign n6310 = n6306 ^ n6300 ;
  assign n6311 = n6310 ^ n6260 ;
  assign n6150 = x119 ^ x115 ;
  assign n6151 = x247 ^ x243 ;
  assign n6163 = n6150 & n6151 ;
  assign n6148 = x118 ^ x114 ;
  assign n6149 = x246 ^ x242 ;
  assign n6162 = n6148 & n6149 ;
  assign n6167 = n6163 ^ n6162 ;
  assign n6146 = x117 ^ x113 ;
  assign n6147 = x245 ^ x241 ;
  assign n6156 = n6146 & n6147 ;
  assign n6144 = x116 ^ x112 ;
  assign n6145 = x244 ^ x240 ;
  assign n6155 = n6144 & n6145 ;
  assign n6160 = n6156 ^ n6155 ;
  assign n6181 = n6167 ^ n6160 ;
  assign n6191 = n6187 ^ n6181 ;
  assign n6192 = n6191 ^ n6141 ;
  assign n6464 = n6311 ^ n6192 ;
  assign n5865 = x111 ^ x107 ;
  assign n5866 = x239 ^ x235 ;
  assign n5878 = n5865 & n5866 ;
  assign n5863 = x110 ^ x106 ;
  assign n5864 = x238 ^ x234 ;
  assign n5877 = n5863 & n5864 ;
  assign n5882 = n5878 ^ n5877 ;
  assign n5861 = x109 ^ x105 ;
  assign n5862 = x237 ^ x233 ;
  assign n5871 = n5861 & n5862 ;
  assign n5859 = x108 ^ x104 ;
  assign n5860 = x236 ^ x232 ;
  assign n5870 = n5859 & n5860 ;
  assign n5875 = n5871 ^ n5870 ;
  assign n5896 = n5882 ^ n5875 ;
  assign n5906 = n5902 ^ n5896 ;
  assign n5907 = n5906 ^ n5856 ;
  assign n5746 = x103 ^ x99 ;
  assign n5747 = x231 ^ x227 ;
  assign n5759 = n5746 & n5747 ;
  assign n5744 = x102 ^ x98 ;
  assign n5745 = x230 ^ x226 ;
  assign n5758 = n5744 & n5745 ;
  assign n5763 = n5759 ^ n5758 ;
  assign n5742 = x101 ^ x97 ;
  assign n5743 = x229 ^ x225 ;
  assign n5752 = n5742 & n5743 ;
  assign n5740 = x100 ^ x96 ;
  assign n5741 = x228 ^ x224 ;
  assign n5751 = n5740 & n5741 ;
  assign n5756 = n5752 ^ n5751 ;
  assign n5777 = n5763 ^ n5756 ;
  assign n5787 = n5783 ^ n5777 ;
  assign n5788 = n5787 ^ n5737 ;
  assign n6060 = n5907 ^ n5788 ;
  assign n6939 = n6464 ^ n6060 ;
  assign n4962 = x95 ^ x91 ;
  assign n4963 = x223 ^ x219 ;
  assign n4975 = n4962 & n4963 ;
  assign n4960 = x94 ^ x90 ;
  assign n4961 = x222 ^ x218 ;
  assign n4974 = n4960 & n4961 ;
  assign n4979 = n4975 ^ n4974 ;
  assign n4958 = x93 ^ x89 ;
  assign n4959 = x221 ^ x217 ;
  assign n4968 = n4958 & n4959 ;
  assign n4956 = x92 ^ x88 ;
  assign n4957 = x220 ^ x216 ;
  assign n4967 = n4956 & n4957 ;
  assign n4972 = n4968 ^ n4967 ;
  assign n4993 = n4979 ^ n4972 ;
  assign n5003 = n4999 ^ n4993 ;
  assign n5004 = n5003 ^ n4953 ;
  assign n4843 = x87 ^ x83 ;
  assign n4844 = x215 ^ x211 ;
  assign n4856 = n4843 & n4844 ;
  assign n4841 = x86 ^ x82 ;
  assign n4842 = x214 ^ x210 ;
  assign n4855 = n4841 & n4842 ;
  assign n4860 = n4856 ^ n4855 ;
  assign n4839 = x85 ^ x81 ;
  assign n4840 = x213 ^ x209 ;
  assign n4849 = n4839 & n4840 ;
  assign n4837 = x84 ^ x80 ;
  assign n4838 = x212 ^ x208 ;
  assign n4848 = n4837 & n4838 ;
  assign n4853 = n4849 ^ n4848 ;
  assign n4874 = n4860 ^ n4853 ;
  assign n4884 = n4880 ^ n4874 ;
  assign n4885 = n4884 ^ n4834 ;
  assign n5157 = n5004 ^ n4885 ;
  assign n4558 = x79 ^ x75 ;
  assign n4559 = x207 ^ x203 ;
  assign n4571 = n4558 & n4559 ;
  assign n4556 = x78 ^ x74 ;
  assign n4557 = x206 ^ x202 ;
  assign n4570 = n4556 & n4557 ;
  assign n4575 = n4571 ^ n4570 ;
  assign n4554 = x77 ^ x73 ;
  assign n4555 = x205 ^ x201 ;
  assign n4564 = n4554 & n4555 ;
  assign n4552 = x76 ^ x72 ;
  assign n4553 = x204 ^ x200 ;
  assign n4563 = n4552 & n4553 ;
  assign n4568 = n4564 ^ n4563 ;
  assign n4589 = n4575 ^ n4568 ;
  assign n4599 = n4595 ^ n4589 ;
  assign n4600 = n4599 ^ n4549 ;
  assign n4439 = x71 ^ x67 ;
  assign n4440 = x199 ^ x195 ;
  assign n4452 = n4439 & n4440 ;
  assign n4437 = x70 ^ x66 ;
  assign n4438 = x198 ^ x194 ;
  assign n4451 = n4437 & n4438 ;
  assign n4456 = n4452 ^ n4451 ;
  assign n4435 = x69 ^ x65 ;
  assign n4436 = x197 ^ x193 ;
  assign n4445 = n4435 & n4436 ;
  assign n4433 = x68 ^ x64 ;
  assign n4434 = x196 ^ x192 ;
  assign n4444 = n4433 & n4434 ;
  assign n4449 = n4445 ^ n4444 ;
  assign n4470 = n4456 ^ n4449 ;
  assign n4480 = n4476 ^ n4470 ;
  assign n4481 = n4480 ^ n4430 ;
  assign n4753 = n4600 ^ n4481 ;
  assign n5632 = n5157 ^ n4753 ;
  assign n8389 = n6939 ^ n5632 ;
  assign n2157 = x63 ^ x59 ;
  assign n2158 = x191 ^ x187 ;
  assign n2170 = n2157 & n2158 ;
  assign n2155 = x62 ^ x58 ;
  assign n2156 = x190 ^ x186 ;
  assign n2169 = n2155 & n2156 ;
  assign n2174 = n2170 ^ n2169 ;
  assign n2153 = x61 ^ x57 ;
  assign n2154 = x189 ^ x185 ;
  assign n2163 = n2153 & n2154 ;
  assign n2151 = x60 ^ x56 ;
  assign n2152 = x188 ^ x184 ;
  assign n2162 = n2151 & n2152 ;
  assign n2167 = n2163 ^ n2162 ;
  assign n2188 = n2174 ^ n2167 ;
  assign n2198 = n2194 ^ n2188 ;
  assign n2199 = n2198 ^ n2148 ;
  assign n2038 = x55 ^ x51 ;
  assign n2039 = x183 ^ x179 ;
  assign n2051 = n2038 & n2039 ;
  assign n2036 = x54 ^ x50 ;
  assign n2037 = x182 ^ x178 ;
  assign n2050 = n2036 & n2037 ;
  assign n2055 = n2051 ^ n2050 ;
  assign n2034 = x53 ^ x49 ;
  assign n2035 = x181 ^ x177 ;
  assign n2044 = n2034 & n2035 ;
  assign n2032 = x52 ^ x48 ;
  assign n2033 = x180 ^ x176 ;
  assign n2043 = n2032 & n2033 ;
  assign n2048 = n2044 ^ n2043 ;
  assign n2069 = n2055 ^ n2048 ;
  assign n2079 = n2075 ^ n2069 ;
  assign n2080 = n2079 ^ n2029 ;
  assign n2352 = n2199 ^ n2080 ;
  assign n1753 = x47 ^ x43 ;
  assign n1754 = x175 ^ x171 ;
  assign n1766 = n1753 & n1754 ;
  assign n1751 = x46 ^ x42 ;
  assign n1752 = x174 ^ x170 ;
  assign n1765 = n1751 & n1752 ;
  assign n1770 = n1766 ^ n1765 ;
  assign n1749 = x45 ^ x41 ;
  assign n1750 = x173 ^ x169 ;
  assign n1759 = n1749 & n1750 ;
  assign n1747 = x44 ^ x40 ;
  assign n1748 = x172 ^ x168 ;
  assign n1758 = n1747 & n1748 ;
  assign n1763 = n1759 ^ n1758 ;
  assign n1784 = n1770 ^ n1763 ;
  assign n1794 = n1790 ^ n1784 ;
  assign n1795 = n1794 ^ n1744 ;
  assign n1634 = x39 ^ x35 ;
  assign n1635 = x167 ^ x163 ;
  assign n1647 = n1634 & n1635 ;
  assign n1632 = x38 ^ x34 ;
  assign n1633 = x166 ^ x162 ;
  assign n1646 = n1632 & n1633 ;
  assign n1651 = n1647 ^ n1646 ;
  assign n1630 = x37 ^ x33 ;
  assign n1631 = x165 ^ x161 ;
  assign n1640 = n1630 & n1631 ;
  assign n1628 = x36 ^ x32 ;
  assign n1629 = x164 ^ x160 ;
  assign n1639 = n1628 & n1629 ;
  assign n1644 = n1640 ^ n1639 ;
  assign n1665 = n1651 ^ n1644 ;
  assign n1675 = n1671 ^ n1665 ;
  assign n1676 = n1675 ^ n1625 ;
  assign n1948 = n1795 ^ n1676 ;
  assign n2827 = n2352 ^ n1948 ;
  assign n850 = x31 ^ x27 ;
  assign n851 = x159 ^ x155 ;
  assign n863 = n850 & n851 ;
  assign n848 = x30 ^ x26 ;
  assign n849 = x158 ^ x154 ;
  assign n862 = n848 & n849 ;
  assign n867 = n863 ^ n862 ;
  assign n846 = x29 ^ x25 ;
  assign n847 = x157 ^ x153 ;
  assign n856 = n846 & n847 ;
  assign n844 = x28 ^ x24 ;
  assign n845 = x156 ^ x152 ;
  assign n855 = n844 & n845 ;
  assign n860 = n856 ^ n855 ;
  assign n881 = n867 ^ n860 ;
  assign n891 = n887 ^ n881 ;
  assign n892 = n891 ^ n841 ;
  assign n731 = x23 ^ x19 ;
  assign n732 = x151 ^ x147 ;
  assign n744 = n731 & n732 ;
  assign n729 = x22 ^ x18 ;
  assign n730 = x150 ^ x146 ;
  assign n743 = n729 & n730 ;
  assign n748 = n744 ^ n743 ;
  assign n727 = x21 ^ x17 ;
  assign n728 = x149 ^ x145 ;
  assign n737 = n727 & n728 ;
  assign n725 = x20 ^ x16 ;
  assign n726 = x148 ^ x144 ;
  assign n736 = n725 & n726 ;
  assign n741 = n737 ^ n736 ;
  assign n762 = n748 ^ n741 ;
  assign n772 = n768 ^ n762 ;
  assign n773 = n772 ^ n722 ;
  assign n1045 = n892 ^ n773 ;
  assign n446 = x15 ^ x11 ;
  assign n447 = x143 ^ x139 ;
  assign n459 = n446 & n447 ;
  assign n444 = x14 ^ x10 ;
  assign n445 = x142 ^ x138 ;
  assign n458 = n444 & n445 ;
  assign n463 = n459 ^ n458 ;
  assign n442 = x13 ^ x9 ;
  assign n443 = x141 ^ x137 ;
  assign n452 = n442 & n443 ;
  assign n440 = x12 ^ x8 ;
  assign n441 = x140 ^ x136 ;
  assign n451 = n440 & n441 ;
  assign n456 = n452 ^ n451 ;
  assign n477 = n463 ^ n456 ;
  assign n487 = n483 ^ n477 ;
  assign n488 = n487 ^ n437 ;
  assign n327 = x7 ^ x3 ;
  assign n328 = x135 ^ x131 ;
  assign n340 = n327 & n328 ;
  assign n325 = x6 ^ x2 ;
  assign n326 = x134 ^ x130 ;
  assign n339 = n325 & n326 ;
  assign n344 = n340 ^ n339 ;
  assign n323 = x5 ^ x1 ;
  assign n324 = x133 ^ x129 ;
  assign n333 = n323 & n324 ;
  assign n321 = x4 ^ x0 ;
  assign n322 = x132 ^ x128 ;
  assign n332 = n321 & n322 ;
  assign n337 = n333 ^ n332 ;
  assign n358 = n344 ^ n337 ;
  assign n368 = n364 ^ n358 ;
  assign n369 = n368 ^ n318 ;
  assign n641 = n488 ^ n369 ;
  assign n1520 = n1045 ^ n641 ;
  assign n4277 = n2827 ^ n1520 ;
  assign n12788 = n8389 ^ n4277 ;
  assign n6283 = n6269 ^ n6267 ;
  assign n6284 = n6270 ^ n6268 ;
  assign n6285 = n6283 & n6284 ;
  assign n6287 = n6285 ^ n6281 ;
  assign n6276 = n6265 ^ n6263 ;
  assign n6277 = n6266 ^ n6264 ;
  assign n6278 = n6276 & n6277 ;
  assign n6280 = n6278 ^ n6274 ;
  assign n6301 = n6287 ^ n6280 ;
  assign n6312 = n6307 ^ n6301 ;
  assign n6313 = n6312 ^ n6262 ;
  assign n6164 = n6150 ^ n6148 ;
  assign n6165 = n6151 ^ n6149 ;
  assign n6166 = n6164 & n6165 ;
  assign n6168 = n6166 ^ n6162 ;
  assign n6157 = n6146 ^ n6144 ;
  assign n6158 = n6147 ^ n6145 ;
  assign n6159 = n6157 & n6158 ;
  assign n6161 = n6159 ^ n6155 ;
  assign n6182 = n6168 ^ n6161 ;
  assign n6193 = n6188 ^ n6182 ;
  assign n6194 = n6193 ^ n6143 ;
  assign n6465 = n6313 ^ n6194 ;
  assign n5879 = n5865 ^ n5863 ;
  assign n5880 = n5866 ^ n5864 ;
  assign n5881 = n5879 & n5880 ;
  assign n5883 = n5881 ^ n5877 ;
  assign n5872 = n5861 ^ n5859 ;
  assign n5873 = n5862 ^ n5860 ;
  assign n5874 = n5872 & n5873 ;
  assign n5876 = n5874 ^ n5870 ;
  assign n5897 = n5883 ^ n5876 ;
  assign n5908 = n5903 ^ n5897 ;
  assign n5909 = n5908 ^ n5858 ;
  assign n5760 = n5746 ^ n5744 ;
  assign n5761 = n5747 ^ n5745 ;
  assign n5762 = n5760 & n5761 ;
  assign n5764 = n5762 ^ n5758 ;
  assign n5753 = n5742 ^ n5740 ;
  assign n5754 = n5743 ^ n5741 ;
  assign n5755 = n5753 & n5754 ;
  assign n5757 = n5755 ^ n5751 ;
  assign n5778 = n5764 ^ n5757 ;
  assign n5789 = n5784 ^ n5778 ;
  assign n5790 = n5789 ^ n5739 ;
  assign n6061 = n5909 ^ n5790 ;
  assign n6940 = n6465 ^ n6061 ;
  assign n4976 = n4962 ^ n4960 ;
  assign n4977 = n4963 ^ n4961 ;
  assign n4978 = n4976 & n4977 ;
  assign n4980 = n4978 ^ n4974 ;
  assign n4969 = n4958 ^ n4956 ;
  assign n4970 = n4959 ^ n4957 ;
  assign n4971 = n4969 & n4970 ;
  assign n4973 = n4971 ^ n4967 ;
  assign n4994 = n4980 ^ n4973 ;
  assign n5005 = n5000 ^ n4994 ;
  assign n5006 = n5005 ^ n4955 ;
  assign n4857 = n4843 ^ n4841 ;
  assign n4858 = n4844 ^ n4842 ;
  assign n4859 = n4857 & n4858 ;
  assign n4861 = n4859 ^ n4855 ;
  assign n4850 = n4839 ^ n4837 ;
  assign n4851 = n4840 ^ n4838 ;
  assign n4852 = n4850 & n4851 ;
  assign n4854 = n4852 ^ n4848 ;
  assign n4875 = n4861 ^ n4854 ;
  assign n4886 = n4881 ^ n4875 ;
  assign n4887 = n4886 ^ n4836 ;
  assign n5158 = n5006 ^ n4887 ;
  assign n4572 = n4558 ^ n4556 ;
  assign n4573 = n4559 ^ n4557 ;
  assign n4574 = n4572 & n4573 ;
  assign n4576 = n4574 ^ n4570 ;
  assign n4565 = n4554 ^ n4552 ;
  assign n4566 = n4555 ^ n4553 ;
  assign n4567 = n4565 & n4566 ;
  assign n4569 = n4567 ^ n4563 ;
  assign n4590 = n4576 ^ n4569 ;
  assign n4601 = n4596 ^ n4590 ;
  assign n4602 = n4601 ^ n4551 ;
  assign n4453 = n4439 ^ n4437 ;
  assign n4454 = n4440 ^ n4438 ;
  assign n4455 = n4453 & n4454 ;
  assign n4457 = n4455 ^ n4451 ;
  assign n4446 = n4435 ^ n4433 ;
  assign n4447 = n4436 ^ n4434 ;
  assign n4448 = n4446 & n4447 ;
  assign n4450 = n4448 ^ n4444 ;
  assign n4471 = n4457 ^ n4450 ;
  assign n4482 = n4477 ^ n4471 ;
  assign n4483 = n4482 ^ n4432 ;
  assign n4754 = n4602 ^ n4483 ;
  assign n5633 = n5158 ^ n4754 ;
  assign n8390 = n6940 ^ n5633 ;
  assign n2171 = n2157 ^ n2155 ;
  assign n2172 = n2158 ^ n2156 ;
  assign n2173 = n2171 & n2172 ;
  assign n2175 = n2173 ^ n2169 ;
  assign n2164 = n2153 ^ n2151 ;
  assign n2165 = n2154 ^ n2152 ;
  assign n2166 = n2164 & n2165 ;
  assign n2168 = n2166 ^ n2162 ;
  assign n2189 = n2175 ^ n2168 ;
  assign n2200 = n2195 ^ n2189 ;
  assign n2201 = n2200 ^ n2150 ;
  assign n2052 = n2038 ^ n2036 ;
  assign n2053 = n2039 ^ n2037 ;
  assign n2054 = n2052 & n2053 ;
  assign n2056 = n2054 ^ n2050 ;
  assign n2045 = n2034 ^ n2032 ;
  assign n2046 = n2035 ^ n2033 ;
  assign n2047 = n2045 & n2046 ;
  assign n2049 = n2047 ^ n2043 ;
  assign n2070 = n2056 ^ n2049 ;
  assign n2081 = n2076 ^ n2070 ;
  assign n2082 = n2081 ^ n2031 ;
  assign n2353 = n2201 ^ n2082 ;
  assign n1767 = n1753 ^ n1751 ;
  assign n1768 = n1754 ^ n1752 ;
  assign n1769 = n1767 & n1768 ;
  assign n1771 = n1769 ^ n1765 ;
  assign n1760 = n1749 ^ n1747 ;
  assign n1761 = n1750 ^ n1748 ;
  assign n1762 = n1760 & n1761 ;
  assign n1764 = n1762 ^ n1758 ;
  assign n1785 = n1771 ^ n1764 ;
  assign n1796 = n1791 ^ n1785 ;
  assign n1797 = n1796 ^ n1746 ;
  assign n1648 = n1634 ^ n1632 ;
  assign n1649 = n1635 ^ n1633 ;
  assign n1650 = n1648 & n1649 ;
  assign n1652 = n1650 ^ n1646 ;
  assign n1641 = n1630 ^ n1628 ;
  assign n1642 = n1631 ^ n1629 ;
  assign n1643 = n1641 & n1642 ;
  assign n1645 = n1643 ^ n1639 ;
  assign n1666 = n1652 ^ n1645 ;
  assign n1677 = n1672 ^ n1666 ;
  assign n1678 = n1677 ^ n1627 ;
  assign n1949 = n1797 ^ n1678 ;
  assign n2828 = n2353 ^ n1949 ;
  assign n864 = n850 ^ n848 ;
  assign n865 = n851 ^ n849 ;
  assign n866 = n864 & n865 ;
  assign n868 = n866 ^ n862 ;
  assign n857 = n846 ^ n844 ;
  assign n858 = n847 ^ n845 ;
  assign n859 = n857 & n858 ;
  assign n861 = n859 ^ n855 ;
  assign n882 = n868 ^ n861 ;
  assign n893 = n888 ^ n882 ;
  assign n894 = n893 ^ n843 ;
  assign n745 = n731 ^ n729 ;
  assign n746 = n732 ^ n730 ;
  assign n747 = n745 & n746 ;
  assign n749 = n747 ^ n743 ;
  assign n738 = n727 ^ n725 ;
  assign n739 = n728 ^ n726 ;
  assign n740 = n738 & n739 ;
  assign n742 = n740 ^ n736 ;
  assign n763 = n749 ^ n742 ;
  assign n774 = n769 ^ n763 ;
  assign n775 = n774 ^ n724 ;
  assign n1046 = n894 ^ n775 ;
  assign n460 = n446 ^ n444 ;
  assign n461 = n447 ^ n445 ;
  assign n462 = n460 & n461 ;
  assign n464 = n462 ^ n458 ;
  assign n453 = n442 ^ n440 ;
  assign n454 = n443 ^ n441 ;
  assign n455 = n453 & n454 ;
  assign n457 = n455 ^ n451 ;
  assign n478 = n464 ^ n457 ;
  assign n489 = n484 ^ n478 ;
  assign n490 = n489 ^ n439 ;
  assign n341 = n327 ^ n325 ;
  assign n342 = n328 ^ n326 ;
  assign n343 = n341 & n342 ;
  assign n345 = n343 ^ n339 ;
  assign n334 = n323 ^ n321 ;
  assign n335 = n324 ^ n322 ;
  assign n336 = n334 & n335 ;
  assign n338 = n336 ^ n332 ;
  assign n359 = n345 ^ n338 ;
  assign n370 = n365 ^ n359 ;
  assign n371 = n370 ^ n320 ;
  assign n642 = n490 ^ n371 ;
  assign n1521 = n1046 ^ n642 ;
  assign n4278 = n2828 ^ n1521 ;
  assign n12789 = n8390 ^ n4278 ;
  assign n6290 = n6269 ^ n6265 ;
  assign n6291 = n6270 ^ n6266 ;
  assign n6294 = n6290 & n6291 ;
  assign n6288 = n6267 ^ n6263 ;
  assign n6289 = n6268 ^ n6264 ;
  assign n6293 = n6288 & n6289 ;
  assign n6298 = n6294 ^ n6293 ;
  assign n6302 = n6300 ^ n6298 ;
  assign n6303 = n6302 ^ n6287 ;
  assign n6314 = n6308 ^ n6303 ;
  assign n6272 = n6262 ^ n6257 ;
  assign n6315 = n6314 ^ n6272 ;
  assign n6171 = n6150 ^ n6146 ;
  assign n6172 = n6151 ^ n6147 ;
  assign n6175 = n6171 & n6172 ;
  assign n6169 = n6148 ^ n6144 ;
  assign n6170 = n6149 ^ n6145 ;
  assign n6174 = n6169 & n6170 ;
  assign n6179 = n6175 ^ n6174 ;
  assign n6183 = n6181 ^ n6179 ;
  assign n6184 = n6183 ^ n6168 ;
  assign n6195 = n6189 ^ n6184 ;
  assign n6153 = n6143 ^ n6138 ;
  assign n6196 = n6195 ^ n6153 ;
  assign n6466 = n6315 ^ n6196 ;
  assign n5886 = n5865 ^ n5861 ;
  assign n5887 = n5866 ^ n5862 ;
  assign n5890 = n5886 & n5887 ;
  assign n5884 = n5863 ^ n5859 ;
  assign n5885 = n5864 ^ n5860 ;
  assign n5889 = n5884 & n5885 ;
  assign n5894 = n5890 ^ n5889 ;
  assign n5898 = n5896 ^ n5894 ;
  assign n5899 = n5898 ^ n5883 ;
  assign n5910 = n5904 ^ n5899 ;
  assign n5868 = n5858 ^ n5853 ;
  assign n5911 = n5910 ^ n5868 ;
  assign n5767 = n5746 ^ n5742 ;
  assign n5768 = n5747 ^ n5743 ;
  assign n5771 = n5767 & n5768 ;
  assign n5765 = n5744 ^ n5740 ;
  assign n5766 = n5745 ^ n5741 ;
  assign n5770 = n5765 & n5766 ;
  assign n5775 = n5771 ^ n5770 ;
  assign n5779 = n5777 ^ n5775 ;
  assign n5780 = n5779 ^ n5764 ;
  assign n5791 = n5785 ^ n5780 ;
  assign n5749 = n5739 ^ n5734 ;
  assign n5792 = n5791 ^ n5749 ;
  assign n6062 = n5911 ^ n5792 ;
  assign n6941 = n6466 ^ n6062 ;
  assign n4983 = n4962 ^ n4958 ;
  assign n4984 = n4963 ^ n4959 ;
  assign n4987 = n4983 & n4984 ;
  assign n4981 = n4960 ^ n4956 ;
  assign n4982 = n4961 ^ n4957 ;
  assign n4986 = n4981 & n4982 ;
  assign n4991 = n4987 ^ n4986 ;
  assign n4995 = n4993 ^ n4991 ;
  assign n4996 = n4995 ^ n4980 ;
  assign n5007 = n5001 ^ n4996 ;
  assign n4965 = n4955 ^ n4950 ;
  assign n5008 = n5007 ^ n4965 ;
  assign n4864 = n4843 ^ n4839 ;
  assign n4865 = n4844 ^ n4840 ;
  assign n4868 = n4864 & n4865 ;
  assign n4862 = n4841 ^ n4837 ;
  assign n4863 = n4842 ^ n4838 ;
  assign n4867 = n4862 & n4863 ;
  assign n4872 = n4868 ^ n4867 ;
  assign n4876 = n4874 ^ n4872 ;
  assign n4877 = n4876 ^ n4861 ;
  assign n4888 = n4882 ^ n4877 ;
  assign n4846 = n4836 ^ n4831 ;
  assign n4889 = n4888 ^ n4846 ;
  assign n5159 = n5008 ^ n4889 ;
  assign n4579 = n4558 ^ n4554 ;
  assign n4580 = n4559 ^ n4555 ;
  assign n4583 = n4579 & n4580 ;
  assign n4577 = n4556 ^ n4552 ;
  assign n4578 = n4557 ^ n4553 ;
  assign n4582 = n4577 & n4578 ;
  assign n4587 = n4583 ^ n4582 ;
  assign n4591 = n4589 ^ n4587 ;
  assign n4592 = n4591 ^ n4576 ;
  assign n4603 = n4597 ^ n4592 ;
  assign n4561 = n4551 ^ n4546 ;
  assign n4604 = n4603 ^ n4561 ;
  assign n4460 = n4439 ^ n4435 ;
  assign n4461 = n4440 ^ n4436 ;
  assign n4464 = n4460 & n4461 ;
  assign n4458 = n4437 ^ n4433 ;
  assign n4459 = n4438 ^ n4434 ;
  assign n4463 = n4458 & n4459 ;
  assign n4468 = n4464 ^ n4463 ;
  assign n4472 = n4470 ^ n4468 ;
  assign n4473 = n4472 ^ n4457 ;
  assign n4484 = n4478 ^ n4473 ;
  assign n4442 = n4432 ^ n4427 ;
  assign n4485 = n4484 ^ n4442 ;
  assign n4755 = n4604 ^ n4485 ;
  assign n5634 = n5159 ^ n4755 ;
  assign n8391 = n6941 ^ n5634 ;
  assign n2178 = n2157 ^ n2153 ;
  assign n2179 = n2158 ^ n2154 ;
  assign n2182 = n2178 & n2179 ;
  assign n2176 = n2155 ^ n2151 ;
  assign n2177 = n2156 ^ n2152 ;
  assign n2181 = n2176 & n2177 ;
  assign n2186 = n2182 ^ n2181 ;
  assign n2190 = n2188 ^ n2186 ;
  assign n2191 = n2190 ^ n2175 ;
  assign n2202 = n2196 ^ n2191 ;
  assign n2160 = n2150 ^ n2145 ;
  assign n2203 = n2202 ^ n2160 ;
  assign n2059 = n2038 ^ n2034 ;
  assign n2060 = n2039 ^ n2035 ;
  assign n2063 = n2059 & n2060 ;
  assign n2057 = n2036 ^ n2032 ;
  assign n2058 = n2037 ^ n2033 ;
  assign n2062 = n2057 & n2058 ;
  assign n2067 = n2063 ^ n2062 ;
  assign n2071 = n2069 ^ n2067 ;
  assign n2072 = n2071 ^ n2056 ;
  assign n2083 = n2077 ^ n2072 ;
  assign n2041 = n2031 ^ n2026 ;
  assign n2084 = n2083 ^ n2041 ;
  assign n2354 = n2203 ^ n2084 ;
  assign n1774 = n1753 ^ n1749 ;
  assign n1775 = n1754 ^ n1750 ;
  assign n1778 = n1774 & n1775 ;
  assign n1772 = n1751 ^ n1747 ;
  assign n1773 = n1752 ^ n1748 ;
  assign n1777 = n1772 & n1773 ;
  assign n1782 = n1778 ^ n1777 ;
  assign n1786 = n1784 ^ n1782 ;
  assign n1787 = n1786 ^ n1771 ;
  assign n1798 = n1792 ^ n1787 ;
  assign n1756 = n1746 ^ n1741 ;
  assign n1799 = n1798 ^ n1756 ;
  assign n1655 = n1634 ^ n1630 ;
  assign n1656 = n1635 ^ n1631 ;
  assign n1659 = n1655 & n1656 ;
  assign n1653 = n1632 ^ n1628 ;
  assign n1654 = n1633 ^ n1629 ;
  assign n1658 = n1653 & n1654 ;
  assign n1663 = n1659 ^ n1658 ;
  assign n1667 = n1665 ^ n1663 ;
  assign n1668 = n1667 ^ n1652 ;
  assign n1679 = n1673 ^ n1668 ;
  assign n1637 = n1627 ^ n1622 ;
  assign n1680 = n1679 ^ n1637 ;
  assign n1950 = n1799 ^ n1680 ;
  assign n2829 = n2354 ^ n1950 ;
  assign n871 = n850 ^ n846 ;
  assign n872 = n851 ^ n847 ;
  assign n875 = n871 & n872 ;
  assign n869 = n848 ^ n844 ;
  assign n870 = n849 ^ n845 ;
  assign n874 = n869 & n870 ;
  assign n879 = n875 ^ n874 ;
  assign n883 = n881 ^ n879 ;
  assign n884 = n883 ^ n868 ;
  assign n895 = n889 ^ n884 ;
  assign n853 = n843 ^ n838 ;
  assign n896 = n895 ^ n853 ;
  assign n752 = n731 ^ n727 ;
  assign n753 = n732 ^ n728 ;
  assign n756 = n752 & n753 ;
  assign n750 = n729 ^ n725 ;
  assign n751 = n730 ^ n726 ;
  assign n755 = n750 & n751 ;
  assign n760 = n756 ^ n755 ;
  assign n764 = n762 ^ n760 ;
  assign n765 = n764 ^ n749 ;
  assign n776 = n770 ^ n765 ;
  assign n734 = n724 ^ n719 ;
  assign n777 = n776 ^ n734 ;
  assign n1047 = n896 ^ n777 ;
  assign n467 = n446 ^ n442 ;
  assign n468 = n447 ^ n443 ;
  assign n471 = n467 & n468 ;
  assign n465 = n444 ^ n440 ;
  assign n466 = n445 ^ n441 ;
  assign n470 = n465 & n466 ;
  assign n475 = n471 ^ n470 ;
  assign n479 = n477 ^ n475 ;
  assign n480 = n479 ^ n464 ;
  assign n491 = n485 ^ n480 ;
  assign n449 = n439 ^ n434 ;
  assign n492 = n491 ^ n449 ;
  assign n348 = n327 ^ n323 ;
  assign n349 = n328 ^ n324 ;
  assign n352 = n348 & n349 ;
  assign n346 = n325 ^ n321 ;
  assign n347 = n326 ^ n322 ;
  assign n351 = n346 & n347 ;
  assign n356 = n352 ^ n351 ;
  assign n360 = n358 ^ n356 ;
  assign n361 = n360 ^ n345 ;
  assign n372 = n366 ^ n361 ;
  assign n330 = n320 ^ n315 ;
  assign n373 = n372 ^ n330 ;
  assign n643 = n492 ^ n373 ;
  assign n1522 = n1047 ^ n643 ;
  assign n4279 = n2829 ^ n1522 ;
  assign n12790 = n8391 ^ n4279 ;
  assign n6295 = n6290 ^ n6288 ;
  assign n6296 = n6291 ^ n6289 ;
  assign n6297 = n6295 & n6296 ;
  assign n6299 = n6297 ^ n6293 ;
  assign n6304 = n6301 ^ n6299 ;
  assign n6292 = n6287 ^ n6286 ;
  assign n6305 = n6304 ^ n6292 ;
  assign n6316 = n6309 ^ n6305 ;
  assign n6271 = n6262 ^ n6260 ;
  assign n6273 = n6271 ^ n6258 ;
  assign n6317 = n6316 ^ n6273 ;
  assign n6176 = n6171 ^ n6169 ;
  assign n6177 = n6172 ^ n6170 ;
  assign n6178 = n6176 & n6177 ;
  assign n6180 = n6178 ^ n6174 ;
  assign n6185 = n6182 ^ n6180 ;
  assign n6173 = n6168 ^ n6167 ;
  assign n6186 = n6185 ^ n6173 ;
  assign n6197 = n6190 ^ n6186 ;
  assign n6152 = n6143 ^ n6141 ;
  assign n6154 = n6152 ^ n6139 ;
  assign n6198 = n6197 ^ n6154 ;
  assign n6467 = n6317 ^ n6198 ;
  assign n5891 = n5886 ^ n5884 ;
  assign n5892 = n5887 ^ n5885 ;
  assign n5893 = n5891 & n5892 ;
  assign n5895 = n5893 ^ n5889 ;
  assign n5900 = n5897 ^ n5895 ;
  assign n5888 = n5883 ^ n5882 ;
  assign n5901 = n5900 ^ n5888 ;
  assign n5912 = n5905 ^ n5901 ;
  assign n5867 = n5858 ^ n5856 ;
  assign n5869 = n5867 ^ n5854 ;
  assign n5913 = n5912 ^ n5869 ;
  assign n5772 = n5767 ^ n5765 ;
  assign n5773 = n5768 ^ n5766 ;
  assign n5774 = n5772 & n5773 ;
  assign n5776 = n5774 ^ n5770 ;
  assign n5781 = n5778 ^ n5776 ;
  assign n5769 = n5764 ^ n5763 ;
  assign n5782 = n5781 ^ n5769 ;
  assign n5793 = n5786 ^ n5782 ;
  assign n5748 = n5739 ^ n5737 ;
  assign n5750 = n5748 ^ n5735 ;
  assign n5794 = n5793 ^ n5750 ;
  assign n6063 = n5913 ^ n5794 ;
  assign n6942 = n6467 ^ n6063 ;
  assign n4988 = n4983 ^ n4981 ;
  assign n4989 = n4984 ^ n4982 ;
  assign n4990 = n4988 & n4989 ;
  assign n4992 = n4990 ^ n4986 ;
  assign n4997 = n4994 ^ n4992 ;
  assign n4985 = n4980 ^ n4979 ;
  assign n4998 = n4997 ^ n4985 ;
  assign n5009 = n5002 ^ n4998 ;
  assign n4964 = n4955 ^ n4953 ;
  assign n4966 = n4964 ^ n4951 ;
  assign n5010 = n5009 ^ n4966 ;
  assign n4869 = n4864 ^ n4862 ;
  assign n4870 = n4865 ^ n4863 ;
  assign n4871 = n4869 & n4870 ;
  assign n4873 = n4871 ^ n4867 ;
  assign n4878 = n4875 ^ n4873 ;
  assign n4866 = n4861 ^ n4860 ;
  assign n4879 = n4878 ^ n4866 ;
  assign n4890 = n4883 ^ n4879 ;
  assign n4845 = n4836 ^ n4834 ;
  assign n4847 = n4845 ^ n4832 ;
  assign n4891 = n4890 ^ n4847 ;
  assign n5160 = n5010 ^ n4891 ;
  assign n4584 = n4579 ^ n4577 ;
  assign n4585 = n4580 ^ n4578 ;
  assign n4586 = n4584 & n4585 ;
  assign n4588 = n4586 ^ n4582 ;
  assign n4593 = n4590 ^ n4588 ;
  assign n4581 = n4576 ^ n4575 ;
  assign n4594 = n4593 ^ n4581 ;
  assign n4605 = n4598 ^ n4594 ;
  assign n4560 = n4551 ^ n4549 ;
  assign n4562 = n4560 ^ n4547 ;
  assign n4606 = n4605 ^ n4562 ;
  assign n4465 = n4460 ^ n4458 ;
  assign n4466 = n4461 ^ n4459 ;
  assign n4467 = n4465 & n4466 ;
  assign n4469 = n4467 ^ n4463 ;
  assign n4474 = n4471 ^ n4469 ;
  assign n4462 = n4457 ^ n4456 ;
  assign n4475 = n4474 ^ n4462 ;
  assign n4486 = n4479 ^ n4475 ;
  assign n4441 = n4432 ^ n4430 ;
  assign n4443 = n4441 ^ n4428 ;
  assign n4487 = n4486 ^ n4443 ;
  assign n4756 = n4606 ^ n4487 ;
  assign n5635 = n5160 ^ n4756 ;
  assign n8392 = n6942 ^ n5635 ;
  assign n2183 = n2178 ^ n2176 ;
  assign n2184 = n2179 ^ n2177 ;
  assign n2185 = n2183 & n2184 ;
  assign n2187 = n2185 ^ n2181 ;
  assign n2192 = n2189 ^ n2187 ;
  assign n2180 = n2175 ^ n2174 ;
  assign n2193 = n2192 ^ n2180 ;
  assign n2204 = n2197 ^ n2193 ;
  assign n2159 = n2150 ^ n2148 ;
  assign n2161 = n2159 ^ n2146 ;
  assign n2205 = n2204 ^ n2161 ;
  assign n2064 = n2059 ^ n2057 ;
  assign n2065 = n2060 ^ n2058 ;
  assign n2066 = n2064 & n2065 ;
  assign n2068 = n2066 ^ n2062 ;
  assign n2073 = n2070 ^ n2068 ;
  assign n2061 = n2056 ^ n2055 ;
  assign n2074 = n2073 ^ n2061 ;
  assign n2085 = n2078 ^ n2074 ;
  assign n2040 = n2031 ^ n2029 ;
  assign n2042 = n2040 ^ n2027 ;
  assign n2086 = n2085 ^ n2042 ;
  assign n2355 = n2205 ^ n2086 ;
  assign n1779 = n1774 ^ n1772 ;
  assign n1780 = n1775 ^ n1773 ;
  assign n1781 = n1779 & n1780 ;
  assign n1783 = n1781 ^ n1777 ;
  assign n1788 = n1785 ^ n1783 ;
  assign n1776 = n1771 ^ n1770 ;
  assign n1789 = n1788 ^ n1776 ;
  assign n1800 = n1793 ^ n1789 ;
  assign n1755 = n1746 ^ n1744 ;
  assign n1757 = n1755 ^ n1742 ;
  assign n1801 = n1800 ^ n1757 ;
  assign n1660 = n1655 ^ n1653 ;
  assign n1661 = n1656 ^ n1654 ;
  assign n1662 = n1660 & n1661 ;
  assign n1664 = n1662 ^ n1658 ;
  assign n1669 = n1666 ^ n1664 ;
  assign n1657 = n1652 ^ n1651 ;
  assign n1670 = n1669 ^ n1657 ;
  assign n1681 = n1674 ^ n1670 ;
  assign n1636 = n1627 ^ n1625 ;
  assign n1638 = n1636 ^ n1623 ;
  assign n1682 = n1681 ^ n1638 ;
  assign n1951 = n1801 ^ n1682 ;
  assign n2830 = n2355 ^ n1951 ;
  assign n876 = n871 ^ n869 ;
  assign n877 = n872 ^ n870 ;
  assign n878 = n876 & n877 ;
  assign n880 = n878 ^ n874 ;
  assign n885 = n882 ^ n880 ;
  assign n873 = n868 ^ n867 ;
  assign n886 = n885 ^ n873 ;
  assign n897 = n890 ^ n886 ;
  assign n852 = n843 ^ n841 ;
  assign n854 = n852 ^ n839 ;
  assign n898 = n897 ^ n854 ;
  assign n757 = n752 ^ n750 ;
  assign n758 = n753 ^ n751 ;
  assign n759 = n757 & n758 ;
  assign n761 = n759 ^ n755 ;
  assign n766 = n763 ^ n761 ;
  assign n754 = n749 ^ n748 ;
  assign n767 = n766 ^ n754 ;
  assign n778 = n771 ^ n767 ;
  assign n733 = n724 ^ n722 ;
  assign n735 = n733 ^ n720 ;
  assign n779 = n778 ^ n735 ;
  assign n1048 = n898 ^ n779 ;
  assign n472 = n467 ^ n465 ;
  assign n473 = n468 ^ n466 ;
  assign n474 = n472 & n473 ;
  assign n476 = n474 ^ n470 ;
  assign n481 = n478 ^ n476 ;
  assign n469 = n464 ^ n463 ;
  assign n482 = n481 ^ n469 ;
  assign n493 = n486 ^ n482 ;
  assign n448 = n439 ^ n437 ;
  assign n450 = n448 ^ n435 ;
  assign n494 = n493 ^ n450 ;
  assign n353 = n348 ^ n346 ;
  assign n354 = n349 ^ n347 ;
  assign n355 = n353 & n354 ;
  assign n357 = n355 ^ n351 ;
  assign n362 = n359 ^ n357 ;
  assign n350 = n345 ^ n344 ;
  assign n363 = n362 ^ n350 ;
  assign n374 = n367 ^ n363 ;
  assign n329 = n320 ^ n318 ;
  assign n331 = n329 ^ n316 ;
  assign n375 = n374 ^ n331 ;
  assign n644 = n494 ^ n375 ;
  assign n1523 = n1048 ^ n644 ;
  assign n4280 = n2830 ^ n1523 ;
  assign n12791 = n8392 ^ n4280 ;
  assign n6332 = x127 ^ x119 ;
  assign n6333 = x255 ^ x247 ;
  assign n6381 = n6332 & n6333 ;
  assign n6330 = x126 ^ x118 ;
  assign n6331 = x254 ^ x246 ;
  assign n6380 = n6330 & n6331 ;
  assign n6385 = n6381 ^ n6380 ;
  assign n6328 = x125 ^ x117 ;
  assign n6329 = x253 ^ x245 ;
  assign n6374 = n6328 & n6329 ;
  assign n6326 = x124 ^ x116 ;
  assign n6327 = x252 ^ x244 ;
  assign n6373 = n6326 & n6327 ;
  assign n6378 = n6374 ^ n6373 ;
  assign n6399 = n6385 ^ n6378 ;
  assign n6324 = x123 ^ x115 ;
  assign n6325 = x251 ^ x243 ;
  assign n6349 = n6324 & n6325 ;
  assign n6322 = x122 ^ x114 ;
  assign n6323 = x250 ^ x242 ;
  assign n6348 = n6322 & n6323 ;
  assign n6353 = n6349 ^ n6348 ;
  assign n6320 = x121 ^ x113 ;
  assign n6321 = x249 ^ x241 ;
  assign n6342 = n6320 & n6321 ;
  assign n6318 = x120 ^ x112 ;
  assign n6319 = x248 ^ x240 ;
  assign n6341 = n6318 & n6319 ;
  assign n6346 = n6342 ^ n6341 ;
  assign n6367 = n6353 ^ n6346 ;
  assign n6448 = n6399 ^ n6367 ;
  assign n6468 = n6460 ^ n6448 ;
  assign n6469 = n6468 ^ n6311 ;
  assign n5928 = x111 ^ x103 ;
  assign n5929 = x239 ^ x231 ;
  assign n5977 = n5928 & n5929 ;
  assign n5926 = x110 ^ x102 ;
  assign n5927 = x238 ^ x230 ;
  assign n5976 = n5926 & n5927 ;
  assign n5981 = n5977 ^ n5976 ;
  assign n5924 = x109 ^ x101 ;
  assign n5925 = x237 ^ x229 ;
  assign n5970 = n5924 & n5925 ;
  assign n5922 = x108 ^ x100 ;
  assign n5923 = x236 ^ x228 ;
  assign n5969 = n5922 & n5923 ;
  assign n5974 = n5970 ^ n5969 ;
  assign n5995 = n5981 ^ n5974 ;
  assign n5920 = x107 ^ x99 ;
  assign n5921 = x235 ^ x227 ;
  assign n5945 = n5920 & n5921 ;
  assign n5918 = x106 ^ x98 ;
  assign n5919 = x234 ^ x226 ;
  assign n5944 = n5918 & n5919 ;
  assign n5949 = n5945 ^ n5944 ;
  assign n5916 = x105 ^ x97 ;
  assign n5917 = x233 ^ x225 ;
  assign n5938 = n5916 & n5917 ;
  assign n5914 = x104 ^ x96 ;
  assign n5915 = x232 ^ x224 ;
  assign n5937 = n5914 & n5915 ;
  assign n5942 = n5938 ^ n5937 ;
  assign n5963 = n5949 ^ n5942 ;
  assign n6044 = n5995 ^ n5963 ;
  assign n6064 = n6056 ^ n6044 ;
  assign n6065 = n6064 ^ n5907 ;
  assign n6943 = n6469 ^ n6065 ;
  assign n5025 = x95 ^ x87 ;
  assign n5026 = x223 ^ x215 ;
  assign n5074 = n5025 & n5026 ;
  assign n5023 = x94 ^ x86 ;
  assign n5024 = x222 ^ x214 ;
  assign n5073 = n5023 & n5024 ;
  assign n5078 = n5074 ^ n5073 ;
  assign n5021 = x93 ^ x85 ;
  assign n5022 = x221 ^ x213 ;
  assign n5067 = n5021 & n5022 ;
  assign n5019 = x92 ^ x84 ;
  assign n5020 = x220 ^ x212 ;
  assign n5066 = n5019 & n5020 ;
  assign n5071 = n5067 ^ n5066 ;
  assign n5092 = n5078 ^ n5071 ;
  assign n5017 = x91 ^ x83 ;
  assign n5018 = x219 ^ x211 ;
  assign n5042 = n5017 & n5018 ;
  assign n5015 = x90 ^ x82 ;
  assign n5016 = x218 ^ x210 ;
  assign n5041 = n5015 & n5016 ;
  assign n5046 = n5042 ^ n5041 ;
  assign n5013 = x89 ^ x81 ;
  assign n5014 = x217 ^ x209 ;
  assign n5035 = n5013 & n5014 ;
  assign n5011 = x88 ^ x80 ;
  assign n5012 = x216 ^ x208 ;
  assign n5034 = n5011 & n5012 ;
  assign n5039 = n5035 ^ n5034 ;
  assign n5060 = n5046 ^ n5039 ;
  assign n5141 = n5092 ^ n5060 ;
  assign n5161 = n5153 ^ n5141 ;
  assign n5162 = n5161 ^ n5004 ;
  assign n4621 = x79 ^ x71 ;
  assign n4622 = x207 ^ x199 ;
  assign n4670 = n4621 & n4622 ;
  assign n4619 = x78 ^ x70 ;
  assign n4620 = x206 ^ x198 ;
  assign n4669 = n4619 & n4620 ;
  assign n4674 = n4670 ^ n4669 ;
  assign n4617 = x77 ^ x69 ;
  assign n4618 = x205 ^ x197 ;
  assign n4663 = n4617 & n4618 ;
  assign n4615 = x76 ^ x68 ;
  assign n4616 = x204 ^ x196 ;
  assign n4662 = n4615 & n4616 ;
  assign n4667 = n4663 ^ n4662 ;
  assign n4688 = n4674 ^ n4667 ;
  assign n4613 = x75 ^ x67 ;
  assign n4614 = x203 ^ x195 ;
  assign n4638 = n4613 & n4614 ;
  assign n4611 = x74 ^ x66 ;
  assign n4612 = x202 ^ x194 ;
  assign n4637 = n4611 & n4612 ;
  assign n4642 = n4638 ^ n4637 ;
  assign n4609 = x73 ^ x65 ;
  assign n4610 = x201 ^ x193 ;
  assign n4631 = n4609 & n4610 ;
  assign n4607 = x72 ^ x64 ;
  assign n4608 = x200 ^ x192 ;
  assign n4630 = n4607 & n4608 ;
  assign n4635 = n4631 ^ n4630 ;
  assign n4656 = n4642 ^ n4635 ;
  assign n4737 = n4688 ^ n4656 ;
  assign n4757 = n4749 ^ n4737 ;
  assign n4758 = n4757 ^ n4600 ;
  assign n5636 = n5162 ^ n4758 ;
  assign n8393 = n6943 ^ n5636 ;
  assign n2220 = x63 ^ x55 ;
  assign n2221 = x191 ^ x183 ;
  assign n2269 = n2220 & n2221 ;
  assign n2218 = x62 ^ x54 ;
  assign n2219 = x190 ^ x182 ;
  assign n2268 = n2218 & n2219 ;
  assign n2273 = n2269 ^ n2268 ;
  assign n2216 = x61 ^ x53 ;
  assign n2217 = x189 ^ x181 ;
  assign n2262 = n2216 & n2217 ;
  assign n2214 = x60 ^ x52 ;
  assign n2215 = x188 ^ x180 ;
  assign n2261 = n2214 & n2215 ;
  assign n2266 = n2262 ^ n2261 ;
  assign n2287 = n2273 ^ n2266 ;
  assign n2212 = x59 ^ x51 ;
  assign n2213 = x187 ^ x179 ;
  assign n2237 = n2212 & n2213 ;
  assign n2210 = x58 ^ x50 ;
  assign n2211 = x186 ^ x178 ;
  assign n2236 = n2210 & n2211 ;
  assign n2241 = n2237 ^ n2236 ;
  assign n2208 = x57 ^ x49 ;
  assign n2209 = x185 ^ x177 ;
  assign n2230 = n2208 & n2209 ;
  assign n2206 = x56 ^ x48 ;
  assign n2207 = x184 ^ x176 ;
  assign n2229 = n2206 & n2207 ;
  assign n2234 = n2230 ^ n2229 ;
  assign n2255 = n2241 ^ n2234 ;
  assign n2336 = n2287 ^ n2255 ;
  assign n2356 = n2348 ^ n2336 ;
  assign n2357 = n2356 ^ n2199 ;
  assign n1816 = x47 ^ x39 ;
  assign n1817 = x175 ^ x167 ;
  assign n1865 = n1816 & n1817 ;
  assign n1814 = x46 ^ x38 ;
  assign n1815 = x174 ^ x166 ;
  assign n1864 = n1814 & n1815 ;
  assign n1869 = n1865 ^ n1864 ;
  assign n1812 = x45 ^ x37 ;
  assign n1813 = x173 ^ x165 ;
  assign n1858 = n1812 & n1813 ;
  assign n1810 = x44 ^ x36 ;
  assign n1811 = x172 ^ x164 ;
  assign n1857 = n1810 & n1811 ;
  assign n1862 = n1858 ^ n1857 ;
  assign n1883 = n1869 ^ n1862 ;
  assign n1808 = x43 ^ x35 ;
  assign n1809 = x171 ^ x163 ;
  assign n1833 = n1808 & n1809 ;
  assign n1806 = x42 ^ x34 ;
  assign n1807 = x170 ^ x162 ;
  assign n1832 = n1806 & n1807 ;
  assign n1837 = n1833 ^ n1832 ;
  assign n1804 = x41 ^ x33 ;
  assign n1805 = x169 ^ x161 ;
  assign n1826 = n1804 & n1805 ;
  assign n1802 = x40 ^ x32 ;
  assign n1803 = x168 ^ x160 ;
  assign n1825 = n1802 & n1803 ;
  assign n1830 = n1826 ^ n1825 ;
  assign n1851 = n1837 ^ n1830 ;
  assign n1932 = n1883 ^ n1851 ;
  assign n1952 = n1944 ^ n1932 ;
  assign n1953 = n1952 ^ n1795 ;
  assign n2831 = n2357 ^ n1953 ;
  assign n913 = x31 ^ x23 ;
  assign n914 = x159 ^ x151 ;
  assign n962 = n913 & n914 ;
  assign n911 = x30 ^ x22 ;
  assign n912 = x158 ^ x150 ;
  assign n961 = n911 & n912 ;
  assign n966 = n962 ^ n961 ;
  assign n909 = x29 ^ x21 ;
  assign n910 = x157 ^ x149 ;
  assign n955 = n909 & n910 ;
  assign n907 = x28 ^ x20 ;
  assign n908 = x156 ^ x148 ;
  assign n954 = n907 & n908 ;
  assign n959 = n955 ^ n954 ;
  assign n980 = n966 ^ n959 ;
  assign n905 = x27 ^ x19 ;
  assign n906 = x155 ^ x147 ;
  assign n930 = n905 & n906 ;
  assign n903 = x26 ^ x18 ;
  assign n904 = x154 ^ x146 ;
  assign n929 = n903 & n904 ;
  assign n934 = n930 ^ n929 ;
  assign n901 = x25 ^ x17 ;
  assign n902 = x153 ^ x145 ;
  assign n923 = n901 & n902 ;
  assign n899 = x24 ^ x16 ;
  assign n900 = x152 ^ x144 ;
  assign n922 = n899 & n900 ;
  assign n927 = n923 ^ n922 ;
  assign n948 = n934 ^ n927 ;
  assign n1029 = n980 ^ n948 ;
  assign n1049 = n1041 ^ n1029 ;
  assign n1050 = n1049 ^ n892 ;
  assign n509 = x15 ^ x7 ;
  assign n510 = x143 ^ x135 ;
  assign n558 = n509 & n510 ;
  assign n507 = x14 ^ x6 ;
  assign n508 = x142 ^ x134 ;
  assign n557 = n507 & n508 ;
  assign n562 = n558 ^ n557 ;
  assign n505 = x13 ^ x5 ;
  assign n506 = x141 ^ x133 ;
  assign n551 = n505 & n506 ;
  assign n503 = x12 ^ x4 ;
  assign n504 = x140 ^ x132 ;
  assign n550 = n503 & n504 ;
  assign n555 = n551 ^ n550 ;
  assign n576 = n562 ^ n555 ;
  assign n501 = x11 ^ x3 ;
  assign n502 = x139 ^ x131 ;
  assign n526 = n501 & n502 ;
  assign n499 = x10 ^ x2 ;
  assign n500 = x138 ^ x130 ;
  assign n525 = n499 & n500 ;
  assign n530 = n526 ^ n525 ;
  assign n497 = x9 ^ x1 ;
  assign n498 = x137 ^ x129 ;
  assign n519 = n497 & n498 ;
  assign n495 = x8 ^ x0 ;
  assign n496 = x136 ^ x128 ;
  assign n518 = n495 & n496 ;
  assign n523 = n519 ^ n518 ;
  assign n544 = n530 ^ n523 ;
  assign n625 = n576 ^ n544 ;
  assign n645 = n637 ^ n625 ;
  assign n646 = n645 ^ n488 ;
  assign n1524 = n1050 ^ n646 ;
  assign n4281 = n2831 ^ n1524 ;
  assign n12792 = n8393 ^ n4281 ;
  assign n6382 = n6332 ^ n6330 ;
  assign n6383 = n6333 ^ n6331 ;
  assign n6384 = n6382 & n6383 ;
  assign n6386 = n6384 ^ n6380 ;
  assign n6375 = n6328 ^ n6326 ;
  assign n6376 = n6329 ^ n6327 ;
  assign n6377 = n6375 & n6376 ;
  assign n6379 = n6377 ^ n6373 ;
  assign n6400 = n6386 ^ n6379 ;
  assign n6350 = n6324 ^ n6322 ;
  assign n6351 = n6325 ^ n6323 ;
  assign n6352 = n6350 & n6351 ;
  assign n6354 = n6352 ^ n6348 ;
  assign n6343 = n6320 ^ n6318 ;
  assign n6344 = n6321 ^ n6319 ;
  assign n6345 = n6343 & n6344 ;
  assign n6347 = n6345 ^ n6341 ;
  assign n6368 = n6354 ^ n6347 ;
  assign n6449 = n6400 ^ n6368 ;
  assign n6470 = n6461 ^ n6449 ;
  assign n6471 = n6470 ^ n6313 ;
  assign n5978 = n5928 ^ n5926 ;
  assign n5979 = n5929 ^ n5927 ;
  assign n5980 = n5978 & n5979 ;
  assign n5982 = n5980 ^ n5976 ;
  assign n5971 = n5924 ^ n5922 ;
  assign n5972 = n5925 ^ n5923 ;
  assign n5973 = n5971 & n5972 ;
  assign n5975 = n5973 ^ n5969 ;
  assign n5996 = n5982 ^ n5975 ;
  assign n5946 = n5920 ^ n5918 ;
  assign n5947 = n5921 ^ n5919 ;
  assign n5948 = n5946 & n5947 ;
  assign n5950 = n5948 ^ n5944 ;
  assign n5939 = n5916 ^ n5914 ;
  assign n5940 = n5917 ^ n5915 ;
  assign n5941 = n5939 & n5940 ;
  assign n5943 = n5941 ^ n5937 ;
  assign n5964 = n5950 ^ n5943 ;
  assign n6045 = n5996 ^ n5964 ;
  assign n6066 = n6057 ^ n6045 ;
  assign n6067 = n6066 ^ n5909 ;
  assign n6944 = n6471 ^ n6067 ;
  assign n5075 = n5025 ^ n5023 ;
  assign n5076 = n5026 ^ n5024 ;
  assign n5077 = n5075 & n5076 ;
  assign n5079 = n5077 ^ n5073 ;
  assign n5068 = n5021 ^ n5019 ;
  assign n5069 = n5022 ^ n5020 ;
  assign n5070 = n5068 & n5069 ;
  assign n5072 = n5070 ^ n5066 ;
  assign n5093 = n5079 ^ n5072 ;
  assign n5043 = n5017 ^ n5015 ;
  assign n5044 = n5018 ^ n5016 ;
  assign n5045 = n5043 & n5044 ;
  assign n5047 = n5045 ^ n5041 ;
  assign n5036 = n5013 ^ n5011 ;
  assign n5037 = n5014 ^ n5012 ;
  assign n5038 = n5036 & n5037 ;
  assign n5040 = n5038 ^ n5034 ;
  assign n5061 = n5047 ^ n5040 ;
  assign n5142 = n5093 ^ n5061 ;
  assign n5163 = n5154 ^ n5142 ;
  assign n5164 = n5163 ^ n5006 ;
  assign n4671 = n4621 ^ n4619 ;
  assign n4672 = n4622 ^ n4620 ;
  assign n4673 = n4671 & n4672 ;
  assign n4675 = n4673 ^ n4669 ;
  assign n4664 = n4617 ^ n4615 ;
  assign n4665 = n4618 ^ n4616 ;
  assign n4666 = n4664 & n4665 ;
  assign n4668 = n4666 ^ n4662 ;
  assign n4689 = n4675 ^ n4668 ;
  assign n4639 = n4613 ^ n4611 ;
  assign n4640 = n4614 ^ n4612 ;
  assign n4641 = n4639 & n4640 ;
  assign n4643 = n4641 ^ n4637 ;
  assign n4632 = n4609 ^ n4607 ;
  assign n4633 = n4610 ^ n4608 ;
  assign n4634 = n4632 & n4633 ;
  assign n4636 = n4634 ^ n4630 ;
  assign n4657 = n4643 ^ n4636 ;
  assign n4738 = n4689 ^ n4657 ;
  assign n4759 = n4750 ^ n4738 ;
  assign n4760 = n4759 ^ n4602 ;
  assign n5637 = n5164 ^ n4760 ;
  assign n8394 = n6944 ^ n5637 ;
  assign n2270 = n2220 ^ n2218 ;
  assign n2271 = n2221 ^ n2219 ;
  assign n2272 = n2270 & n2271 ;
  assign n2274 = n2272 ^ n2268 ;
  assign n2263 = n2216 ^ n2214 ;
  assign n2264 = n2217 ^ n2215 ;
  assign n2265 = n2263 & n2264 ;
  assign n2267 = n2265 ^ n2261 ;
  assign n2288 = n2274 ^ n2267 ;
  assign n2238 = n2212 ^ n2210 ;
  assign n2239 = n2213 ^ n2211 ;
  assign n2240 = n2238 & n2239 ;
  assign n2242 = n2240 ^ n2236 ;
  assign n2231 = n2208 ^ n2206 ;
  assign n2232 = n2209 ^ n2207 ;
  assign n2233 = n2231 & n2232 ;
  assign n2235 = n2233 ^ n2229 ;
  assign n2256 = n2242 ^ n2235 ;
  assign n2337 = n2288 ^ n2256 ;
  assign n2358 = n2349 ^ n2337 ;
  assign n2359 = n2358 ^ n2201 ;
  assign n1866 = n1816 ^ n1814 ;
  assign n1867 = n1817 ^ n1815 ;
  assign n1868 = n1866 & n1867 ;
  assign n1870 = n1868 ^ n1864 ;
  assign n1859 = n1812 ^ n1810 ;
  assign n1860 = n1813 ^ n1811 ;
  assign n1861 = n1859 & n1860 ;
  assign n1863 = n1861 ^ n1857 ;
  assign n1884 = n1870 ^ n1863 ;
  assign n1834 = n1808 ^ n1806 ;
  assign n1835 = n1809 ^ n1807 ;
  assign n1836 = n1834 & n1835 ;
  assign n1838 = n1836 ^ n1832 ;
  assign n1827 = n1804 ^ n1802 ;
  assign n1828 = n1805 ^ n1803 ;
  assign n1829 = n1827 & n1828 ;
  assign n1831 = n1829 ^ n1825 ;
  assign n1852 = n1838 ^ n1831 ;
  assign n1933 = n1884 ^ n1852 ;
  assign n1954 = n1945 ^ n1933 ;
  assign n1955 = n1954 ^ n1797 ;
  assign n2832 = n2359 ^ n1955 ;
  assign n963 = n913 ^ n911 ;
  assign n964 = n914 ^ n912 ;
  assign n965 = n963 & n964 ;
  assign n967 = n965 ^ n961 ;
  assign n956 = n909 ^ n907 ;
  assign n957 = n910 ^ n908 ;
  assign n958 = n956 & n957 ;
  assign n960 = n958 ^ n954 ;
  assign n981 = n967 ^ n960 ;
  assign n931 = n905 ^ n903 ;
  assign n932 = n906 ^ n904 ;
  assign n933 = n931 & n932 ;
  assign n935 = n933 ^ n929 ;
  assign n924 = n901 ^ n899 ;
  assign n925 = n902 ^ n900 ;
  assign n926 = n924 & n925 ;
  assign n928 = n926 ^ n922 ;
  assign n949 = n935 ^ n928 ;
  assign n1030 = n981 ^ n949 ;
  assign n1051 = n1042 ^ n1030 ;
  assign n1052 = n1051 ^ n894 ;
  assign n559 = n509 ^ n507 ;
  assign n560 = n510 ^ n508 ;
  assign n561 = n559 & n560 ;
  assign n563 = n561 ^ n557 ;
  assign n552 = n505 ^ n503 ;
  assign n553 = n506 ^ n504 ;
  assign n554 = n552 & n553 ;
  assign n556 = n554 ^ n550 ;
  assign n577 = n563 ^ n556 ;
  assign n527 = n501 ^ n499 ;
  assign n528 = n502 ^ n500 ;
  assign n529 = n527 & n528 ;
  assign n531 = n529 ^ n525 ;
  assign n520 = n497 ^ n495 ;
  assign n521 = n498 ^ n496 ;
  assign n522 = n520 & n521 ;
  assign n524 = n522 ^ n518 ;
  assign n545 = n531 ^ n524 ;
  assign n626 = n577 ^ n545 ;
  assign n647 = n638 ^ n626 ;
  assign n648 = n647 ^ n490 ;
  assign n1525 = n1052 ^ n648 ;
  assign n4282 = n2832 ^ n1525 ;
  assign n12793 = n8394 ^ n4282 ;
  assign n6389 = n6332 ^ n6328 ;
  assign n6390 = n6333 ^ n6329 ;
  assign n6393 = n6389 & n6390 ;
  assign n6387 = n6330 ^ n6326 ;
  assign n6388 = n6331 ^ n6327 ;
  assign n6392 = n6387 & n6388 ;
  assign n6397 = n6393 ^ n6392 ;
  assign n6401 = n6399 ^ n6397 ;
  assign n6402 = n6401 ^ n6386 ;
  assign n6357 = n6324 ^ n6320 ;
  assign n6358 = n6325 ^ n6321 ;
  assign n6361 = n6357 & n6358 ;
  assign n6355 = n6322 ^ n6318 ;
  assign n6356 = n6323 ^ n6319 ;
  assign n6360 = n6355 & n6356 ;
  assign n6365 = n6361 ^ n6360 ;
  assign n6369 = n6367 ^ n6365 ;
  assign n6370 = n6369 ^ n6354 ;
  assign n6450 = n6402 ^ n6370 ;
  assign n6472 = n6462 ^ n6450 ;
  assign n6473 = n6472 ^ n6315 ;
  assign n5985 = n5928 ^ n5924 ;
  assign n5986 = n5929 ^ n5925 ;
  assign n5989 = n5985 & n5986 ;
  assign n5983 = n5926 ^ n5922 ;
  assign n5984 = n5927 ^ n5923 ;
  assign n5988 = n5983 & n5984 ;
  assign n5993 = n5989 ^ n5988 ;
  assign n5997 = n5995 ^ n5993 ;
  assign n5998 = n5997 ^ n5982 ;
  assign n5953 = n5920 ^ n5916 ;
  assign n5954 = n5921 ^ n5917 ;
  assign n5957 = n5953 & n5954 ;
  assign n5951 = n5918 ^ n5914 ;
  assign n5952 = n5919 ^ n5915 ;
  assign n5956 = n5951 & n5952 ;
  assign n5961 = n5957 ^ n5956 ;
  assign n5965 = n5963 ^ n5961 ;
  assign n5966 = n5965 ^ n5950 ;
  assign n6046 = n5998 ^ n5966 ;
  assign n6068 = n6058 ^ n6046 ;
  assign n6069 = n6068 ^ n5911 ;
  assign n6945 = n6473 ^ n6069 ;
  assign n5082 = n5025 ^ n5021 ;
  assign n5083 = n5026 ^ n5022 ;
  assign n5086 = n5082 & n5083 ;
  assign n5080 = n5023 ^ n5019 ;
  assign n5081 = n5024 ^ n5020 ;
  assign n5085 = n5080 & n5081 ;
  assign n5090 = n5086 ^ n5085 ;
  assign n5094 = n5092 ^ n5090 ;
  assign n5095 = n5094 ^ n5079 ;
  assign n5050 = n5017 ^ n5013 ;
  assign n5051 = n5018 ^ n5014 ;
  assign n5054 = n5050 & n5051 ;
  assign n5048 = n5015 ^ n5011 ;
  assign n5049 = n5016 ^ n5012 ;
  assign n5053 = n5048 & n5049 ;
  assign n5058 = n5054 ^ n5053 ;
  assign n5062 = n5060 ^ n5058 ;
  assign n5063 = n5062 ^ n5047 ;
  assign n5143 = n5095 ^ n5063 ;
  assign n5165 = n5155 ^ n5143 ;
  assign n5166 = n5165 ^ n5008 ;
  assign n4678 = n4621 ^ n4617 ;
  assign n4679 = n4622 ^ n4618 ;
  assign n4682 = n4678 & n4679 ;
  assign n4676 = n4619 ^ n4615 ;
  assign n4677 = n4620 ^ n4616 ;
  assign n4681 = n4676 & n4677 ;
  assign n4686 = n4682 ^ n4681 ;
  assign n4690 = n4688 ^ n4686 ;
  assign n4691 = n4690 ^ n4675 ;
  assign n4646 = n4613 ^ n4609 ;
  assign n4647 = n4614 ^ n4610 ;
  assign n4650 = n4646 & n4647 ;
  assign n4644 = n4611 ^ n4607 ;
  assign n4645 = n4612 ^ n4608 ;
  assign n4649 = n4644 & n4645 ;
  assign n4654 = n4650 ^ n4649 ;
  assign n4658 = n4656 ^ n4654 ;
  assign n4659 = n4658 ^ n4643 ;
  assign n4739 = n4691 ^ n4659 ;
  assign n4761 = n4751 ^ n4739 ;
  assign n4762 = n4761 ^ n4604 ;
  assign n5638 = n5166 ^ n4762 ;
  assign n8395 = n6945 ^ n5638 ;
  assign n2277 = n2220 ^ n2216 ;
  assign n2278 = n2221 ^ n2217 ;
  assign n2281 = n2277 & n2278 ;
  assign n2275 = n2218 ^ n2214 ;
  assign n2276 = n2219 ^ n2215 ;
  assign n2280 = n2275 & n2276 ;
  assign n2285 = n2281 ^ n2280 ;
  assign n2289 = n2287 ^ n2285 ;
  assign n2290 = n2289 ^ n2274 ;
  assign n2245 = n2212 ^ n2208 ;
  assign n2246 = n2213 ^ n2209 ;
  assign n2249 = n2245 & n2246 ;
  assign n2243 = n2210 ^ n2206 ;
  assign n2244 = n2211 ^ n2207 ;
  assign n2248 = n2243 & n2244 ;
  assign n2253 = n2249 ^ n2248 ;
  assign n2257 = n2255 ^ n2253 ;
  assign n2258 = n2257 ^ n2242 ;
  assign n2338 = n2290 ^ n2258 ;
  assign n2360 = n2350 ^ n2338 ;
  assign n2361 = n2360 ^ n2203 ;
  assign n1873 = n1816 ^ n1812 ;
  assign n1874 = n1817 ^ n1813 ;
  assign n1877 = n1873 & n1874 ;
  assign n1871 = n1814 ^ n1810 ;
  assign n1872 = n1815 ^ n1811 ;
  assign n1876 = n1871 & n1872 ;
  assign n1881 = n1877 ^ n1876 ;
  assign n1885 = n1883 ^ n1881 ;
  assign n1886 = n1885 ^ n1870 ;
  assign n1841 = n1808 ^ n1804 ;
  assign n1842 = n1809 ^ n1805 ;
  assign n1845 = n1841 & n1842 ;
  assign n1839 = n1806 ^ n1802 ;
  assign n1840 = n1807 ^ n1803 ;
  assign n1844 = n1839 & n1840 ;
  assign n1849 = n1845 ^ n1844 ;
  assign n1853 = n1851 ^ n1849 ;
  assign n1854 = n1853 ^ n1838 ;
  assign n1934 = n1886 ^ n1854 ;
  assign n1956 = n1946 ^ n1934 ;
  assign n1957 = n1956 ^ n1799 ;
  assign n2833 = n2361 ^ n1957 ;
  assign n970 = n913 ^ n909 ;
  assign n971 = n914 ^ n910 ;
  assign n974 = n970 & n971 ;
  assign n968 = n911 ^ n907 ;
  assign n969 = n912 ^ n908 ;
  assign n973 = n968 & n969 ;
  assign n978 = n974 ^ n973 ;
  assign n982 = n980 ^ n978 ;
  assign n983 = n982 ^ n967 ;
  assign n938 = n905 ^ n901 ;
  assign n939 = n906 ^ n902 ;
  assign n942 = n938 & n939 ;
  assign n936 = n903 ^ n899 ;
  assign n937 = n904 ^ n900 ;
  assign n941 = n936 & n937 ;
  assign n946 = n942 ^ n941 ;
  assign n950 = n948 ^ n946 ;
  assign n951 = n950 ^ n935 ;
  assign n1031 = n983 ^ n951 ;
  assign n1053 = n1043 ^ n1031 ;
  assign n1054 = n1053 ^ n896 ;
  assign n566 = n509 ^ n505 ;
  assign n567 = n510 ^ n506 ;
  assign n570 = n566 & n567 ;
  assign n564 = n507 ^ n503 ;
  assign n565 = n508 ^ n504 ;
  assign n569 = n564 & n565 ;
  assign n574 = n570 ^ n569 ;
  assign n578 = n576 ^ n574 ;
  assign n579 = n578 ^ n563 ;
  assign n534 = n501 ^ n497 ;
  assign n535 = n502 ^ n498 ;
  assign n538 = n534 & n535 ;
  assign n532 = n499 ^ n495 ;
  assign n533 = n500 ^ n496 ;
  assign n537 = n532 & n533 ;
  assign n542 = n538 ^ n537 ;
  assign n546 = n544 ^ n542 ;
  assign n547 = n546 ^ n531 ;
  assign n627 = n579 ^ n547 ;
  assign n649 = n639 ^ n627 ;
  assign n650 = n649 ^ n492 ;
  assign n1526 = n1054 ^ n650 ;
  assign n4283 = n2833 ^ n1526 ;
  assign n12794 = n8395 ^ n4283 ;
  assign n6394 = n6389 ^ n6387 ;
  assign n6395 = n6390 ^ n6388 ;
  assign n6396 = n6394 & n6395 ;
  assign n6398 = n6396 ^ n6392 ;
  assign n6403 = n6400 ^ n6398 ;
  assign n6391 = n6386 ^ n6385 ;
  assign n6404 = n6403 ^ n6391 ;
  assign n6362 = n6357 ^ n6355 ;
  assign n6363 = n6358 ^ n6356 ;
  assign n6364 = n6362 & n6363 ;
  assign n6366 = n6364 ^ n6360 ;
  assign n6371 = n6368 ^ n6366 ;
  assign n6359 = n6354 ^ n6353 ;
  assign n6372 = n6371 ^ n6359 ;
  assign n6451 = n6404 ^ n6372 ;
  assign n6474 = n6463 ^ n6451 ;
  assign n6475 = n6474 ^ n6317 ;
  assign n5990 = n5985 ^ n5983 ;
  assign n5991 = n5986 ^ n5984 ;
  assign n5992 = n5990 & n5991 ;
  assign n5994 = n5992 ^ n5988 ;
  assign n5999 = n5996 ^ n5994 ;
  assign n5987 = n5982 ^ n5981 ;
  assign n6000 = n5999 ^ n5987 ;
  assign n5958 = n5953 ^ n5951 ;
  assign n5959 = n5954 ^ n5952 ;
  assign n5960 = n5958 & n5959 ;
  assign n5962 = n5960 ^ n5956 ;
  assign n5967 = n5964 ^ n5962 ;
  assign n5955 = n5950 ^ n5949 ;
  assign n5968 = n5967 ^ n5955 ;
  assign n6047 = n6000 ^ n5968 ;
  assign n6070 = n6059 ^ n6047 ;
  assign n6071 = n6070 ^ n5913 ;
  assign n6946 = n6475 ^ n6071 ;
  assign n5087 = n5082 ^ n5080 ;
  assign n5088 = n5083 ^ n5081 ;
  assign n5089 = n5087 & n5088 ;
  assign n5091 = n5089 ^ n5085 ;
  assign n5096 = n5093 ^ n5091 ;
  assign n5084 = n5079 ^ n5078 ;
  assign n5097 = n5096 ^ n5084 ;
  assign n5055 = n5050 ^ n5048 ;
  assign n5056 = n5051 ^ n5049 ;
  assign n5057 = n5055 & n5056 ;
  assign n5059 = n5057 ^ n5053 ;
  assign n5064 = n5061 ^ n5059 ;
  assign n5052 = n5047 ^ n5046 ;
  assign n5065 = n5064 ^ n5052 ;
  assign n5144 = n5097 ^ n5065 ;
  assign n5167 = n5156 ^ n5144 ;
  assign n5168 = n5167 ^ n5010 ;
  assign n4683 = n4678 ^ n4676 ;
  assign n4684 = n4679 ^ n4677 ;
  assign n4685 = n4683 & n4684 ;
  assign n4687 = n4685 ^ n4681 ;
  assign n4692 = n4689 ^ n4687 ;
  assign n4680 = n4675 ^ n4674 ;
  assign n4693 = n4692 ^ n4680 ;
  assign n4651 = n4646 ^ n4644 ;
  assign n4652 = n4647 ^ n4645 ;
  assign n4653 = n4651 & n4652 ;
  assign n4655 = n4653 ^ n4649 ;
  assign n4660 = n4657 ^ n4655 ;
  assign n4648 = n4643 ^ n4642 ;
  assign n4661 = n4660 ^ n4648 ;
  assign n4740 = n4693 ^ n4661 ;
  assign n4763 = n4752 ^ n4740 ;
  assign n4764 = n4763 ^ n4606 ;
  assign n5639 = n5168 ^ n4764 ;
  assign n8396 = n6946 ^ n5639 ;
  assign n2282 = n2277 ^ n2275 ;
  assign n2283 = n2278 ^ n2276 ;
  assign n2284 = n2282 & n2283 ;
  assign n2286 = n2284 ^ n2280 ;
  assign n2291 = n2288 ^ n2286 ;
  assign n2279 = n2274 ^ n2273 ;
  assign n2292 = n2291 ^ n2279 ;
  assign n2250 = n2245 ^ n2243 ;
  assign n2251 = n2246 ^ n2244 ;
  assign n2252 = n2250 & n2251 ;
  assign n2254 = n2252 ^ n2248 ;
  assign n2259 = n2256 ^ n2254 ;
  assign n2247 = n2242 ^ n2241 ;
  assign n2260 = n2259 ^ n2247 ;
  assign n2339 = n2292 ^ n2260 ;
  assign n2362 = n2351 ^ n2339 ;
  assign n2363 = n2362 ^ n2205 ;
  assign n1878 = n1873 ^ n1871 ;
  assign n1879 = n1874 ^ n1872 ;
  assign n1880 = n1878 & n1879 ;
  assign n1882 = n1880 ^ n1876 ;
  assign n1887 = n1884 ^ n1882 ;
  assign n1875 = n1870 ^ n1869 ;
  assign n1888 = n1887 ^ n1875 ;
  assign n1846 = n1841 ^ n1839 ;
  assign n1847 = n1842 ^ n1840 ;
  assign n1848 = n1846 & n1847 ;
  assign n1850 = n1848 ^ n1844 ;
  assign n1855 = n1852 ^ n1850 ;
  assign n1843 = n1838 ^ n1837 ;
  assign n1856 = n1855 ^ n1843 ;
  assign n1935 = n1888 ^ n1856 ;
  assign n1958 = n1947 ^ n1935 ;
  assign n1959 = n1958 ^ n1801 ;
  assign n2834 = n2363 ^ n1959 ;
  assign n975 = n970 ^ n968 ;
  assign n976 = n971 ^ n969 ;
  assign n977 = n975 & n976 ;
  assign n979 = n977 ^ n973 ;
  assign n984 = n981 ^ n979 ;
  assign n972 = n967 ^ n966 ;
  assign n985 = n984 ^ n972 ;
  assign n943 = n938 ^ n936 ;
  assign n944 = n939 ^ n937 ;
  assign n945 = n943 & n944 ;
  assign n947 = n945 ^ n941 ;
  assign n952 = n949 ^ n947 ;
  assign n940 = n935 ^ n934 ;
  assign n953 = n952 ^ n940 ;
  assign n1032 = n985 ^ n953 ;
  assign n1055 = n1044 ^ n1032 ;
  assign n1056 = n1055 ^ n898 ;
  assign n571 = n566 ^ n564 ;
  assign n572 = n567 ^ n565 ;
  assign n573 = n571 & n572 ;
  assign n575 = n573 ^ n569 ;
  assign n580 = n577 ^ n575 ;
  assign n568 = n563 ^ n562 ;
  assign n581 = n580 ^ n568 ;
  assign n539 = n534 ^ n532 ;
  assign n540 = n535 ^ n533 ;
  assign n541 = n539 & n540 ;
  assign n543 = n541 ^ n537 ;
  assign n548 = n545 ^ n543 ;
  assign n536 = n531 ^ n530 ;
  assign n549 = n548 ^ n536 ;
  assign n628 = n581 ^ n549 ;
  assign n651 = n640 ^ n628 ;
  assign n652 = n651 ^ n494 ;
  assign n1527 = n1056 ^ n652 ;
  assign n4284 = n2834 ^ n1527 ;
  assign n12795 = n8396 ^ n4284 ;
  assign n6411 = n6332 ^ n6324 ;
  assign n6412 = n6333 ^ n6325 ;
  assign n6424 = n6411 & n6412 ;
  assign n6409 = n6330 ^ n6322 ;
  assign n6410 = n6331 ^ n6323 ;
  assign n6423 = n6409 & n6410 ;
  assign n6428 = n6424 ^ n6423 ;
  assign n6407 = n6328 ^ n6320 ;
  assign n6408 = n6329 ^ n6321 ;
  assign n6417 = n6407 & n6408 ;
  assign n6405 = n6326 ^ n6318 ;
  assign n6406 = n6327 ^ n6319 ;
  assign n6416 = n6405 & n6406 ;
  assign n6421 = n6417 ^ n6416 ;
  assign n6442 = n6428 ^ n6421 ;
  assign n6452 = n6448 ^ n6442 ;
  assign n6453 = n6452 ^ n6402 ;
  assign n6476 = n6464 ^ n6453 ;
  assign n6337 = n6315 ^ n6306 ;
  assign n6477 = n6476 ^ n6337 ;
  assign n6007 = n5928 ^ n5920 ;
  assign n6008 = n5929 ^ n5921 ;
  assign n6020 = n6007 & n6008 ;
  assign n6005 = n5926 ^ n5918 ;
  assign n6006 = n5927 ^ n5919 ;
  assign n6019 = n6005 & n6006 ;
  assign n6024 = n6020 ^ n6019 ;
  assign n6003 = n5924 ^ n5916 ;
  assign n6004 = n5925 ^ n5917 ;
  assign n6013 = n6003 & n6004 ;
  assign n6001 = n5922 ^ n5914 ;
  assign n6002 = n5923 ^ n5915 ;
  assign n6012 = n6001 & n6002 ;
  assign n6017 = n6013 ^ n6012 ;
  assign n6038 = n6024 ^ n6017 ;
  assign n6048 = n6044 ^ n6038 ;
  assign n6049 = n6048 ^ n5998 ;
  assign n6072 = n6060 ^ n6049 ;
  assign n5933 = n5911 ^ n5902 ;
  assign n6073 = n6072 ^ n5933 ;
  assign n6947 = n6477 ^ n6073 ;
  assign n5104 = n5025 ^ n5017 ;
  assign n5105 = n5026 ^ n5018 ;
  assign n5117 = n5104 & n5105 ;
  assign n5102 = n5023 ^ n5015 ;
  assign n5103 = n5024 ^ n5016 ;
  assign n5116 = n5102 & n5103 ;
  assign n5121 = n5117 ^ n5116 ;
  assign n5100 = n5021 ^ n5013 ;
  assign n5101 = n5022 ^ n5014 ;
  assign n5110 = n5100 & n5101 ;
  assign n5098 = n5019 ^ n5011 ;
  assign n5099 = n5020 ^ n5012 ;
  assign n5109 = n5098 & n5099 ;
  assign n5114 = n5110 ^ n5109 ;
  assign n5135 = n5121 ^ n5114 ;
  assign n5145 = n5141 ^ n5135 ;
  assign n5146 = n5145 ^ n5095 ;
  assign n5169 = n5157 ^ n5146 ;
  assign n5030 = n5008 ^ n4999 ;
  assign n5170 = n5169 ^ n5030 ;
  assign n4700 = n4621 ^ n4613 ;
  assign n4701 = n4622 ^ n4614 ;
  assign n4713 = n4700 & n4701 ;
  assign n4698 = n4619 ^ n4611 ;
  assign n4699 = n4620 ^ n4612 ;
  assign n4712 = n4698 & n4699 ;
  assign n4717 = n4713 ^ n4712 ;
  assign n4696 = n4617 ^ n4609 ;
  assign n4697 = n4618 ^ n4610 ;
  assign n4706 = n4696 & n4697 ;
  assign n4694 = n4615 ^ n4607 ;
  assign n4695 = n4616 ^ n4608 ;
  assign n4705 = n4694 & n4695 ;
  assign n4710 = n4706 ^ n4705 ;
  assign n4731 = n4717 ^ n4710 ;
  assign n4741 = n4737 ^ n4731 ;
  assign n4742 = n4741 ^ n4691 ;
  assign n4765 = n4753 ^ n4742 ;
  assign n4626 = n4604 ^ n4595 ;
  assign n4766 = n4765 ^ n4626 ;
  assign n5640 = n5170 ^ n4766 ;
  assign n8397 = n6947 ^ n5640 ;
  assign n2299 = n2220 ^ n2212 ;
  assign n2300 = n2221 ^ n2213 ;
  assign n2312 = n2299 & n2300 ;
  assign n2297 = n2218 ^ n2210 ;
  assign n2298 = n2219 ^ n2211 ;
  assign n2311 = n2297 & n2298 ;
  assign n2316 = n2312 ^ n2311 ;
  assign n2295 = n2216 ^ n2208 ;
  assign n2296 = n2217 ^ n2209 ;
  assign n2305 = n2295 & n2296 ;
  assign n2293 = n2214 ^ n2206 ;
  assign n2294 = n2215 ^ n2207 ;
  assign n2304 = n2293 & n2294 ;
  assign n2309 = n2305 ^ n2304 ;
  assign n2330 = n2316 ^ n2309 ;
  assign n2340 = n2336 ^ n2330 ;
  assign n2341 = n2340 ^ n2290 ;
  assign n2364 = n2352 ^ n2341 ;
  assign n2225 = n2203 ^ n2194 ;
  assign n2365 = n2364 ^ n2225 ;
  assign n1895 = n1816 ^ n1808 ;
  assign n1896 = n1817 ^ n1809 ;
  assign n1908 = n1895 & n1896 ;
  assign n1893 = n1814 ^ n1806 ;
  assign n1894 = n1815 ^ n1807 ;
  assign n1907 = n1893 & n1894 ;
  assign n1912 = n1908 ^ n1907 ;
  assign n1891 = n1812 ^ n1804 ;
  assign n1892 = n1813 ^ n1805 ;
  assign n1901 = n1891 & n1892 ;
  assign n1889 = n1810 ^ n1802 ;
  assign n1890 = n1811 ^ n1803 ;
  assign n1900 = n1889 & n1890 ;
  assign n1905 = n1901 ^ n1900 ;
  assign n1926 = n1912 ^ n1905 ;
  assign n1936 = n1932 ^ n1926 ;
  assign n1937 = n1936 ^ n1886 ;
  assign n1960 = n1948 ^ n1937 ;
  assign n1821 = n1799 ^ n1790 ;
  assign n1961 = n1960 ^ n1821 ;
  assign n2835 = n2365 ^ n1961 ;
  assign n992 = n913 ^ n905 ;
  assign n993 = n914 ^ n906 ;
  assign n1005 = n992 & n993 ;
  assign n990 = n911 ^ n903 ;
  assign n991 = n912 ^ n904 ;
  assign n1004 = n990 & n991 ;
  assign n1009 = n1005 ^ n1004 ;
  assign n988 = n909 ^ n901 ;
  assign n989 = n910 ^ n902 ;
  assign n998 = n988 & n989 ;
  assign n986 = n907 ^ n899 ;
  assign n987 = n908 ^ n900 ;
  assign n997 = n986 & n987 ;
  assign n1002 = n998 ^ n997 ;
  assign n1023 = n1009 ^ n1002 ;
  assign n1033 = n1029 ^ n1023 ;
  assign n1034 = n1033 ^ n983 ;
  assign n1057 = n1045 ^ n1034 ;
  assign n918 = n896 ^ n887 ;
  assign n1058 = n1057 ^ n918 ;
  assign n588 = n509 ^ n501 ;
  assign n589 = n510 ^ n502 ;
  assign n601 = n588 & n589 ;
  assign n586 = n507 ^ n499 ;
  assign n587 = n508 ^ n500 ;
  assign n600 = n586 & n587 ;
  assign n605 = n601 ^ n600 ;
  assign n584 = n505 ^ n497 ;
  assign n585 = n506 ^ n498 ;
  assign n594 = n584 & n585 ;
  assign n582 = n503 ^ n495 ;
  assign n583 = n504 ^ n496 ;
  assign n593 = n582 & n583 ;
  assign n598 = n594 ^ n593 ;
  assign n619 = n605 ^ n598 ;
  assign n629 = n625 ^ n619 ;
  assign n630 = n629 ^ n579 ;
  assign n653 = n641 ^ n630 ;
  assign n514 = n492 ^ n483 ;
  assign n654 = n653 ^ n514 ;
  assign n1528 = n1058 ^ n654 ;
  assign n4285 = n2835 ^ n1528 ;
  assign n12796 = n8397 ^ n4285 ;
  assign n6425 = n6411 ^ n6409 ;
  assign n6426 = n6412 ^ n6410 ;
  assign n6427 = n6425 & n6426 ;
  assign n6429 = n6427 ^ n6423 ;
  assign n6418 = n6407 ^ n6405 ;
  assign n6419 = n6408 ^ n6406 ;
  assign n6420 = n6418 & n6419 ;
  assign n6422 = n6420 ^ n6416 ;
  assign n6443 = n6429 ^ n6422 ;
  assign n6454 = n6449 ^ n6443 ;
  assign n6455 = n6454 ^ n6404 ;
  assign n6478 = n6465 ^ n6455 ;
  assign n6338 = n6317 ^ n6307 ;
  assign n6479 = n6478 ^ n6338 ;
  assign n6021 = n6007 ^ n6005 ;
  assign n6022 = n6008 ^ n6006 ;
  assign n6023 = n6021 & n6022 ;
  assign n6025 = n6023 ^ n6019 ;
  assign n6014 = n6003 ^ n6001 ;
  assign n6015 = n6004 ^ n6002 ;
  assign n6016 = n6014 & n6015 ;
  assign n6018 = n6016 ^ n6012 ;
  assign n6039 = n6025 ^ n6018 ;
  assign n6050 = n6045 ^ n6039 ;
  assign n6051 = n6050 ^ n6000 ;
  assign n6074 = n6061 ^ n6051 ;
  assign n5934 = n5913 ^ n5903 ;
  assign n6075 = n6074 ^ n5934 ;
  assign n6948 = n6479 ^ n6075 ;
  assign n5118 = n5104 ^ n5102 ;
  assign n5119 = n5105 ^ n5103 ;
  assign n5120 = n5118 & n5119 ;
  assign n5122 = n5120 ^ n5116 ;
  assign n5111 = n5100 ^ n5098 ;
  assign n5112 = n5101 ^ n5099 ;
  assign n5113 = n5111 & n5112 ;
  assign n5115 = n5113 ^ n5109 ;
  assign n5136 = n5122 ^ n5115 ;
  assign n5147 = n5142 ^ n5136 ;
  assign n5148 = n5147 ^ n5097 ;
  assign n5171 = n5158 ^ n5148 ;
  assign n5031 = n5010 ^ n5000 ;
  assign n5172 = n5171 ^ n5031 ;
  assign n4714 = n4700 ^ n4698 ;
  assign n4715 = n4701 ^ n4699 ;
  assign n4716 = n4714 & n4715 ;
  assign n4718 = n4716 ^ n4712 ;
  assign n4707 = n4696 ^ n4694 ;
  assign n4708 = n4697 ^ n4695 ;
  assign n4709 = n4707 & n4708 ;
  assign n4711 = n4709 ^ n4705 ;
  assign n4732 = n4718 ^ n4711 ;
  assign n4743 = n4738 ^ n4732 ;
  assign n4744 = n4743 ^ n4693 ;
  assign n4767 = n4754 ^ n4744 ;
  assign n4627 = n4606 ^ n4596 ;
  assign n4768 = n4767 ^ n4627 ;
  assign n5641 = n5172 ^ n4768 ;
  assign n8398 = n6948 ^ n5641 ;
  assign n2313 = n2299 ^ n2297 ;
  assign n2314 = n2300 ^ n2298 ;
  assign n2315 = n2313 & n2314 ;
  assign n2317 = n2315 ^ n2311 ;
  assign n2306 = n2295 ^ n2293 ;
  assign n2307 = n2296 ^ n2294 ;
  assign n2308 = n2306 & n2307 ;
  assign n2310 = n2308 ^ n2304 ;
  assign n2331 = n2317 ^ n2310 ;
  assign n2342 = n2337 ^ n2331 ;
  assign n2343 = n2342 ^ n2292 ;
  assign n2366 = n2353 ^ n2343 ;
  assign n2226 = n2205 ^ n2195 ;
  assign n2367 = n2366 ^ n2226 ;
  assign n1909 = n1895 ^ n1893 ;
  assign n1910 = n1896 ^ n1894 ;
  assign n1911 = n1909 & n1910 ;
  assign n1913 = n1911 ^ n1907 ;
  assign n1902 = n1891 ^ n1889 ;
  assign n1903 = n1892 ^ n1890 ;
  assign n1904 = n1902 & n1903 ;
  assign n1906 = n1904 ^ n1900 ;
  assign n1927 = n1913 ^ n1906 ;
  assign n1938 = n1933 ^ n1927 ;
  assign n1939 = n1938 ^ n1888 ;
  assign n1962 = n1949 ^ n1939 ;
  assign n1822 = n1801 ^ n1791 ;
  assign n1963 = n1962 ^ n1822 ;
  assign n2836 = n2367 ^ n1963 ;
  assign n1006 = n992 ^ n990 ;
  assign n1007 = n993 ^ n991 ;
  assign n1008 = n1006 & n1007 ;
  assign n1010 = n1008 ^ n1004 ;
  assign n999 = n988 ^ n986 ;
  assign n1000 = n989 ^ n987 ;
  assign n1001 = n999 & n1000 ;
  assign n1003 = n1001 ^ n997 ;
  assign n1024 = n1010 ^ n1003 ;
  assign n1035 = n1030 ^ n1024 ;
  assign n1036 = n1035 ^ n985 ;
  assign n1059 = n1046 ^ n1036 ;
  assign n919 = n898 ^ n888 ;
  assign n1060 = n1059 ^ n919 ;
  assign n602 = n588 ^ n586 ;
  assign n603 = n589 ^ n587 ;
  assign n604 = n602 & n603 ;
  assign n606 = n604 ^ n600 ;
  assign n595 = n584 ^ n582 ;
  assign n596 = n585 ^ n583 ;
  assign n597 = n595 & n596 ;
  assign n599 = n597 ^ n593 ;
  assign n620 = n606 ^ n599 ;
  assign n631 = n626 ^ n620 ;
  assign n632 = n631 ^ n581 ;
  assign n655 = n642 ^ n632 ;
  assign n515 = n494 ^ n484 ;
  assign n656 = n655 ^ n515 ;
  assign n1529 = n1060 ^ n656 ;
  assign n4286 = n2836 ^ n1529 ;
  assign n12797 = n8398 ^ n4286 ;
  assign n6432 = n6411 ^ n6407 ;
  assign n6433 = n6412 ^ n6408 ;
  assign n6436 = n6432 & n6433 ;
  assign n6430 = n6409 ^ n6405 ;
  assign n6431 = n6410 ^ n6406 ;
  assign n6435 = n6430 & n6431 ;
  assign n6440 = n6436 ^ n6435 ;
  assign n6444 = n6442 ^ n6440 ;
  assign n6445 = n6444 ^ n6429 ;
  assign n6456 = n6450 ^ n6445 ;
  assign n6414 = n6404 ^ n6399 ;
  assign n6457 = n6456 ^ n6414 ;
  assign n6480 = n6466 ^ n6457 ;
  assign n6335 = n6317 ^ n6311 ;
  assign n6339 = n6335 ^ n6308 ;
  assign n6481 = n6480 ^ n6339 ;
  assign n6028 = n6007 ^ n6003 ;
  assign n6029 = n6008 ^ n6004 ;
  assign n6032 = n6028 & n6029 ;
  assign n6026 = n6005 ^ n6001 ;
  assign n6027 = n6006 ^ n6002 ;
  assign n6031 = n6026 & n6027 ;
  assign n6036 = n6032 ^ n6031 ;
  assign n6040 = n6038 ^ n6036 ;
  assign n6041 = n6040 ^ n6025 ;
  assign n6052 = n6046 ^ n6041 ;
  assign n6010 = n6000 ^ n5995 ;
  assign n6053 = n6052 ^ n6010 ;
  assign n6076 = n6062 ^ n6053 ;
  assign n5931 = n5913 ^ n5907 ;
  assign n5935 = n5931 ^ n5904 ;
  assign n6077 = n6076 ^ n5935 ;
  assign n6949 = n6481 ^ n6077 ;
  assign n5125 = n5104 ^ n5100 ;
  assign n5126 = n5105 ^ n5101 ;
  assign n5129 = n5125 & n5126 ;
  assign n5123 = n5102 ^ n5098 ;
  assign n5124 = n5103 ^ n5099 ;
  assign n5128 = n5123 & n5124 ;
  assign n5133 = n5129 ^ n5128 ;
  assign n5137 = n5135 ^ n5133 ;
  assign n5138 = n5137 ^ n5122 ;
  assign n5149 = n5143 ^ n5138 ;
  assign n5107 = n5097 ^ n5092 ;
  assign n5150 = n5149 ^ n5107 ;
  assign n5173 = n5159 ^ n5150 ;
  assign n5028 = n5010 ^ n5004 ;
  assign n5032 = n5028 ^ n5001 ;
  assign n5174 = n5173 ^ n5032 ;
  assign n4721 = n4700 ^ n4696 ;
  assign n4722 = n4701 ^ n4697 ;
  assign n4725 = n4721 & n4722 ;
  assign n4719 = n4698 ^ n4694 ;
  assign n4720 = n4699 ^ n4695 ;
  assign n4724 = n4719 & n4720 ;
  assign n4729 = n4725 ^ n4724 ;
  assign n4733 = n4731 ^ n4729 ;
  assign n4734 = n4733 ^ n4718 ;
  assign n4745 = n4739 ^ n4734 ;
  assign n4703 = n4693 ^ n4688 ;
  assign n4746 = n4745 ^ n4703 ;
  assign n4769 = n4755 ^ n4746 ;
  assign n4624 = n4606 ^ n4600 ;
  assign n4628 = n4624 ^ n4597 ;
  assign n4770 = n4769 ^ n4628 ;
  assign n5642 = n5174 ^ n4770 ;
  assign n8399 = n6949 ^ n5642 ;
  assign n2320 = n2299 ^ n2295 ;
  assign n2321 = n2300 ^ n2296 ;
  assign n2324 = n2320 & n2321 ;
  assign n2318 = n2297 ^ n2293 ;
  assign n2319 = n2298 ^ n2294 ;
  assign n2323 = n2318 & n2319 ;
  assign n2328 = n2324 ^ n2323 ;
  assign n2332 = n2330 ^ n2328 ;
  assign n2333 = n2332 ^ n2317 ;
  assign n2344 = n2338 ^ n2333 ;
  assign n2302 = n2292 ^ n2287 ;
  assign n2345 = n2344 ^ n2302 ;
  assign n2368 = n2354 ^ n2345 ;
  assign n2223 = n2205 ^ n2199 ;
  assign n2227 = n2223 ^ n2196 ;
  assign n2369 = n2368 ^ n2227 ;
  assign n1916 = n1895 ^ n1891 ;
  assign n1917 = n1896 ^ n1892 ;
  assign n1920 = n1916 & n1917 ;
  assign n1914 = n1893 ^ n1889 ;
  assign n1915 = n1894 ^ n1890 ;
  assign n1919 = n1914 & n1915 ;
  assign n1924 = n1920 ^ n1919 ;
  assign n1928 = n1926 ^ n1924 ;
  assign n1929 = n1928 ^ n1913 ;
  assign n1940 = n1934 ^ n1929 ;
  assign n1898 = n1888 ^ n1883 ;
  assign n1941 = n1940 ^ n1898 ;
  assign n1964 = n1950 ^ n1941 ;
  assign n1819 = n1801 ^ n1795 ;
  assign n1823 = n1819 ^ n1792 ;
  assign n1965 = n1964 ^ n1823 ;
  assign n2837 = n2369 ^ n1965 ;
  assign n1013 = n992 ^ n988 ;
  assign n1014 = n993 ^ n989 ;
  assign n1017 = n1013 & n1014 ;
  assign n1011 = n990 ^ n986 ;
  assign n1012 = n991 ^ n987 ;
  assign n1016 = n1011 & n1012 ;
  assign n1021 = n1017 ^ n1016 ;
  assign n1025 = n1023 ^ n1021 ;
  assign n1026 = n1025 ^ n1010 ;
  assign n1037 = n1031 ^ n1026 ;
  assign n995 = n985 ^ n980 ;
  assign n1038 = n1037 ^ n995 ;
  assign n1061 = n1047 ^ n1038 ;
  assign n916 = n898 ^ n892 ;
  assign n920 = n916 ^ n889 ;
  assign n1062 = n1061 ^ n920 ;
  assign n609 = n588 ^ n584 ;
  assign n610 = n589 ^ n585 ;
  assign n613 = n609 & n610 ;
  assign n607 = n586 ^ n582 ;
  assign n608 = n587 ^ n583 ;
  assign n612 = n607 & n608 ;
  assign n617 = n613 ^ n612 ;
  assign n621 = n619 ^ n617 ;
  assign n622 = n621 ^ n606 ;
  assign n633 = n627 ^ n622 ;
  assign n591 = n581 ^ n576 ;
  assign n634 = n633 ^ n591 ;
  assign n657 = n643 ^ n634 ;
  assign n512 = n494 ^ n488 ;
  assign n516 = n512 ^ n485 ;
  assign n658 = n657 ^ n516 ;
  assign n1530 = n1062 ^ n658 ;
  assign n4287 = n2837 ^ n1530 ;
  assign n12798 = n8399 ^ n4287 ;
  assign n6437 = n6432 ^ n6430 ;
  assign n6438 = n6433 ^ n6431 ;
  assign n6439 = n6437 & n6438 ;
  assign n6441 = n6439 ^ n6435 ;
  assign n6446 = n6443 ^ n6441 ;
  assign n6434 = n6429 ^ n6428 ;
  assign n6447 = n6446 ^ n6434 ;
  assign n6458 = n6451 ^ n6447 ;
  assign n6413 = n6404 ^ n6402 ;
  assign n6415 = n6413 ^ n6400 ;
  assign n6459 = n6458 ^ n6415 ;
  assign n6482 = n6467 ^ n6459 ;
  assign n6334 = n6317 ^ n6315 ;
  assign n6336 = n6334 ^ n6313 ;
  assign n6340 = n6336 ^ n6309 ;
  assign n6483 = n6482 ^ n6340 ;
  assign n6033 = n6028 ^ n6026 ;
  assign n6034 = n6029 ^ n6027 ;
  assign n6035 = n6033 & n6034 ;
  assign n6037 = n6035 ^ n6031 ;
  assign n6042 = n6039 ^ n6037 ;
  assign n6030 = n6025 ^ n6024 ;
  assign n6043 = n6042 ^ n6030 ;
  assign n6054 = n6047 ^ n6043 ;
  assign n6009 = n6000 ^ n5998 ;
  assign n6011 = n6009 ^ n5996 ;
  assign n6055 = n6054 ^ n6011 ;
  assign n6078 = n6063 ^ n6055 ;
  assign n5930 = n5913 ^ n5911 ;
  assign n5932 = n5930 ^ n5909 ;
  assign n5936 = n5932 ^ n5905 ;
  assign n6079 = n6078 ^ n5936 ;
  assign n6950 = n6483 ^ n6079 ;
  assign n5130 = n5125 ^ n5123 ;
  assign n5131 = n5126 ^ n5124 ;
  assign n5132 = n5130 & n5131 ;
  assign n5134 = n5132 ^ n5128 ;
  assign n5139 = n5136 ^ n5134 ;
  assign n5127 = n5122 ^ n5121 ;
  assign n5140 = n5139 ^ n5127 ;
  assign n5151 = n5144 ^ n5140 ;
  assign n5106 = n5097 ^ n5095 ;
  assign n5108 = n5106 ^ n5093 ;
  assign n5152 = n5151 ^ n5108 ;
  assign n5175 = n5160 ^ n5152 ;
  assign n5027 = n5010 ^ n5008 ;
  assign n5029 = n5027 ^ n5006 ;
  assign n5033 = n5029 ^ n5002 ;
  assign n5176 = n5175 ^ n5033 ;
  assign n4726 = n4721 ^ n4719 ;
  assign n4727 = n4722 ^ n4720 ;
  assign n4728 = n4726 & n4727 ;
  assign n4730 = n4728 ^ n4724 ;
  assign n4735 = n4732 ^ n4730 ;
  assign n4723 = n4718 ^ n4717 ;
  assign n4736 = n4735 ^ n4723 ;
  assign n4747 = n4740 ^ n4736 ;
  assign n4702 = n4693 ^ n4691 ;
  assign n4704 = n4702 ^ n4689 ;
  assign n4748 = n4747 ^ n4704 ;
  assign n4771 = n4756 ^ n4748 ;
  assign n4623 = n4606 ^ n4604 ;
  assign n4625 = n4623 ^ n4602 ;
  assign n4629 = n4625 ^ n4598 ;
  assign n4772 = n4771 ^ n4629 ;
  assign n5643 = n5176 ^ n4772 ;
  assign n8400 = n6950 ^ n5643 ;
  assign n2325 = n2320 ^ n2318 ;
  assign n2326 = n2321 ^ n2319 ;
  assign n2327 = n2325 & n2326 ;
  assign n2329 = n2327 ^ n2323 ;
  assign n2334 = n2331 ^ n2329 ;
  assign n2322 = n2317 ^ n2316 ;
  assign n2335 = n2334 ^ n2322 ;
  assign n2346 = n2339 ^ n2335 ;
  assign n2301 = n2292 ^ n2290 ;
  assign n2303 = n2301 ^ n2288 ;
  assign n2347 = n2346 ^ n2303 ;
  assign n2370 = n2355 ^ n2347 ;
  assign n2222 = n2205 ^ n2203 ;
  assign n2224 = n2222 ^ n2201 ;
  assign n2228 = n2224 ^ n2197 ;
  assign n2371 = n2370 ^ n2228 ;
  assign n1921 = n1916 ^ n1914 ;
  assign n1922 = n1917 ^ n1915 ;
  assign n1923 = n1921 & n1922 ;
  assign n1925 = n1923 ^ n1919 ;
  assign n1930 = n1927 ^ n1925 ;
  assign n1918 = n1913 ^ n1912 ;
  assign n1931 = n1930 ^ n1918 ;
  assign n1942 = n1935 ^ n1931 ;
  assign n1897 = n1888 ^ n1886 ;
  assign n1899 = n1897 ^ n1884 ;
  assign n1943 = n1942 ^ n1899 ;
  assign n1966 = n1951 ^ n1943 ;
  assign n1818 = n1801 ^ n1799 ;
  assign n1820 = n1818 ^ n1797 ;
  assign n1824 = n1820 ^ n1793 ;
  assign n1967 = n1966 ^ n1824 ;
  assign n2838 = n2371 ^ n1967 ;
  assign n1018 = n1013 ^ n1011 ;
  assign n1019 = n1014 ^ n1012 ;
  assign n1020 = n1018 & n1019 ;
  assign n1022 = n1020 ^ n1016 ;
  assign n1027 = n1024 ^ n1022 ;
  assign n1015 = n1010 ^ n1009 ;
  assign n1028 = n1027 ^ n1015 ;
  assign n1039 = n1032 ^ n1028 ;
  assign n994 = n985 ^ n983 ;
  assign n996 = n994 ^ n981 ;
  assign n1040 = n1039 ^ n996 ;
  assign n1063 = n1048 ^ n1040 ;
  assign n915 = n898 ^ n896 ;
  assign n917 = n915 ^ n894 ;
  assign n921 = n917 ^ n890 ;
  assign n1064 = n1063 ^ n921 ;
  assign n614 = n609 ^ n607 ;
  assign n615 = n610 ^ n608 ;
  assign n616 = n614 & n615 ;
  assign n618 = n616 ^ n612 ;
  assign n623 = n620 ^ n618 ;
  assign n611 = n606 ^ n605 ;
  assign n624 = n623 ^ n611 ;
  assign n635 = n628 ^ n624 ;
  assign n590 = n581 ^ n579 ;
  assign n592 = n590 ^ n577 ;
  assign n636 = n635 ^ n592 ;
  assign n659 = n644 ^ n636 ;
  assign n511 = n494 ^ n492 ;
  assign n513 = n511 ^ n490 ;
  assign n517 = n513 ^ n486 ;
  assign n660 = n659 ^ n517 ;
  assign n1531 = n1064 ^ n660 ;
  assign n4288 = n2838 ^ n1531 ;
  assign n12799 = n8400 ^ n4288 ;
  assign n6514 = x127 ^ x111 ;
  assign n6515 = x255 ^ x239 ;
  assign n6690 = n6514 & n6515 ;
  assign n6512 = x126 ^ x110 ;
  assign n6513 = x254 ^ x238 ;
  assign n6689 = n6512 & n6513 ;
  assign n6694 = n6690 ^ n6689 ;
  assign n6510 = x125 ^ x109 ;
  assign n6511 = x253 ^ x237 ;
  assign n6683 = n6510 & n6511 ;
  assign n6508 = x124 ^ x108 ;
  assign n6509 = x252 ^ x236 ;
  assign n6682 = n6508 & n6509 ;
  assign n6687 = n6683 ^ n6682 ;
  assign n6708 = n6694 ^ n6687 ;
  assign n6506 = x123 ^ x107 ;
  assign n6507 = x251 ^ x235 ;
  assign n6658 = n6506 & n6507 ;
  assign n6504 = x122 ^ x106 ;
  assign n6505 = x250 ^ x234 ;
  assign n6657 = n6504 & n6505 ;
  assign n6662 = n6658 ^ n6657 ;
  assign n6502 = x121 ^ x105 ;
  assign n6503 = x249 ^ x233 ;
  assign n6651 = n6502 & n6503 ;
  assign n6500 = x120 ^ x104 ;
  assign n6501 = x248 ^ x232 ;
  assign n6650 = n6500 & n6501 ;
  assign n6655 = n6651 ^ n6650 ;
  assign n6676 = n6662 ^ n6655 ;
  assign n6757 = n6708 ^ n6676 ;
  assign n6498 = x119 ^ x103 ;
  assign n6499 = x247 ^ x231 ;
  assign n6571 = n6498 & n6499 ;
  assign n6496 = x118 ^ x102 ;
  assign n6497 = x246 ^ x230 ;
  assign n6570 = n6496 & n6497 ;
  assign n6575 = n6571 ^ n6570 ;
  assign n6494 = x117 ^ x101 ;
  assign n6495 = x245 ^ x229 ;
  assign n6564 = n6494 & n6495 ;
  assign n6492 = x116 ^ x100 ;
  assign n6493 = x244 ^ x228 ;
  assign n6563 = n6492 & n6493 ;
  assign n6568 = n6564 ^ n6563 ;
  assign n6589 = n6575 ^ n6568 ;
  assign n6490 = x115 ^ x99 ;
  assign n6491 = x243 ^ x227 ;
  assign n6539 = n6490 & n6491 ;
  assign n6488 = x114 ^ x98 ;
  assign n6489 = x242 ^ x226 ;
  assign n6538 = n6488 & n6489 ;
  assign n6543 = n6539 ^ n6538 ;
  assign n6486 = x113 ^ x97 ;
  assign n6487 = x241 ^ x225 ;
  assign n6532 = n6486 & n6487 ;
  assign n6484 = x112 ^ x96 ;
  assign n6485 = x240 ^ x224 ;
  assign n6531 = n6484 & n6485 ;
  assign n6536 = n6532 ^ n6531 ;
  assign n6557 = n6543 ^ n6536 ;
  assign n6638 = n6589 ^ n6557 ;
  assign n6911 = n6757 ^ n6638 ;
  assign n6951 = n6935 ^ n6911 ;
  assign n6952 = n6951 ^ n6469 ;
  assign n5207 = x95 ^ x79 ;
  assign n5208 = x223 ^ x207 ;
  assign n5383 = n5207 & n5208 ;
  assign n5205 = x94 ^ x78 ;
  assign n5206 = x222 ^ x206 ;
  assign n5382 = n5205 & n5206 ;
  assign n5387 = n5383 ^ n5382 ;
  assign n5203 = x93 ^ x77 ;
  assign n5204 = x221 ^ x205 ;
  assign n5376 = n5203 & n5204 ;
  assign n5201 = x92 ^ x76 ;
  assign n5202 = x220 ^ x204 ;
  assign n5375 = n5201 & n5202 ;
  assign n5380 = n5376 ^ n5375 ;
  assign n5401 = n5387 ^ n5380 ;
  assign n5199 = x91 ^ x75 ;
  assign n5200 = x219 ^ x203 ;
  assign n5351 = n5199 & n5200 ;
  assign n5197 = x90 ^ x74 ;
  assign n5198 = x218 ^ x202 ;
  assign n5350 = n5197 & n5198 ;
  assign n5355 = n5351 ^ n5350 ;
  assign n5195 = x89 ^ x73 ;
  assign n5196 = x217 ^ x201 ;
  assign n5344 = n5195 & n5196 ;
  assign n5193 = x88 ^ x72 ;
  assign n5194 = x216 ^ x200 ;
  assign n5343 = n5193 & n5194 ;
  assign n5348 = n5344 ^ n5343 ;
  assign n5369 = n5355 ^ n5348 ;
  assign n5450 = n5401 ^ n5369 ;
  assign n5191 = x87 ^ x71 ;
  assign n5192 = x215 ^ x199 ;
  assign n5264 = n5191 & n5192 ;
  assign n5189 = x86 ^ x70 ;
  assign n5190 = x214 ^ x198 ;
  assign n5263 = n5189 & n5190 ;
  assign n5268 = n5264 ^ n5263 ;
  assign n5187 = x85 ^ x69 ;
  assign n5188 = x213 ^ x197 ;
  assign n5257 = n5187 & n5188 ;
  assign n5185 = x84 ^ x68 ;
  assign n5186 = x212 ^ x196 ;
  assign n5256 = n5185 & n5186 ;
  assign n5261 = n5257 ^ n5256 ;
  assign n5282 = n5268 ^ n5261 ;
  assign n5183 = x83 ^ x67 ;
  assign n5184 = x211 ^ x195 ;
  assign n5232 = n5183 & n5184 ;
  assign n5181 = x82 ^ x66 ;
  assign n5182 = x210 ^ x194 ;
  assign n5231 = n5181 & n5182 ;
  assign n5236 = n5232 ^ n5231 ;
  assign n5179 = x81 ^ x65 ;
  assign n5180 = x209 ^ x193 ;
  assign n5225 = n5179 & n5180 ;
  assign n5177 = x80 ^ x64 ;
  assign n5178 = x208 ^ x192 ;
  assign n5224 = n5177 & n5178 ;
  assign n5229 = n5225 ^ n5224 ;
  assign n5250 = n5236 ^ n5229 ;
  assign n5331 = n5282 ^ n5250 ;
  assign n5604 = n5450 ^ n5331 ;
  assign n5644 = n5628 ^ n5604 ;
  assign n5645 = n5644 ^ n5162 ;
  assign n8401 = n6952 ^ n5645 ;
  assign n2402 = x63 ^ x47 ;
  assign n2403 = x191 ^ x175 ;
  assign n2578 = n2402 & n2403 ;
  assign n2400 = x62 ^ x46 ;
  assign n2401 = x190 ^ x174 ;
  assign n2577 = n2400 & n2401 ;
  assign n2582 = n2578 ^ n2577 ;
  assign n2398 = x61 ^ x45 ;
  assign n2399 = x189 ^ x173 ;
  assign n2571 = n2398 & n2399 ;
  assign n2396 = x60 ^ x44 ;
  assign n2397 = x188 ^ x172 ;
  assign n2570 = n2396 & n2397 ;
  assign n2575 = n2571 ^ n2570 ;
  assign n2596 = n2582 ^ n2575 ;
  assign n2394 = x59 ^ x43 ;
  assign n2395 = x187 ^ x171 ;
  assign n2546 = n2394 & n2395 ;
  assign n2392 = x58 ^ x42 ;
  assign n2393 = x186 ^ x170 ;
  assign n2545 = n2392 & n2393 ;
  assign n2550 = n2546 ^ n2545 ;
  assign n2390 = x57 ^ x41 ;
  assign n2391 = x185 ^ x169 ;
  assign n2539 = n2390 & n2391 ;
  assign n2388 = x56 ^ x40 ;
  assign n2389 = x184 ^ x168 ;
  assign n2538 = n2388 & n2389 ;
  assign n2543 = n2539 ^ n2538 ;
  assign n2564 = n2550 ^ n2543 ;
  assign n2645 = n2596 ^ n2564 ;
  assign n2386 = x55 ^ x39 ;
  assign n2387 = x183 ^ x167 ;
  assign n2459 = n2386 & n2387 ;
  assign n2384 = x54 ^ x38 ;
  assign n2385 = x182 ^ x166 ;
  assign n2458 = n2384 & n2385 ;
  assign n2463 = n2459 ^ n2458 ;
  assign n2382 = x53 ^ x37 ;
  assign n2383 = x181 ^ x165 ;
  assign n2452 = n2382 & n2383 ;
  assign n2380 = x52 ^ x36 ;
  assign n2381 = x180 ^ x164 ;
  assign n2451 = n2380 & n2381 ;
  assign n2456 = n2452 ^ n2451 ;
  assign n2477 = n2463 ^ n2456 ;
  assign n2378 = x51 ^ x35 ;
  assign n2379 = x179 ^ x163 ;
  assign n2427 = n2378 & n2379 ;
  assign n2376 = x50 ^ x34 ;
  assign n2377 = x178 ^ x162 ;
  assign n2426 = n2376 & n2377 ;
  assign n2431 = n2427 ^ n2426 ;
  assign n2374 = x49 ^ x33 ;
  assign n2375 = x177 ^ x161 ;
  assign n2420 = n2374 & n2375 ;
  assign n2372 = x48 ^ x32 ;
  assign n2373 = x176 ^ x160 ;
  assign n2419 = n2372 & n2373 ;
  assign n2424 = n2420 ^ n2419 ;
  assign n2445 = n2431 ^ n2424 ;
  assign n2526 = n2477 ^ n2445 ;
  assign n2799 = n2645 ^ n2526 ;
  assign n2839 = n2823 ^ n2799 ;
  assign n2840 = n2839 ^ n2357 ;
  assign n1095 = x31 ^ x15 ;
  assign n1096 = x159 ^ x143 ;
  assign n1271 = n1095 & n1096 ;
  assign n1093 = x30 ^ x14 ;
  assign n1094 = x158 ^ x142 ;
  assign n1270 = n1093 & n1094 ;
  assign n1275 = n1271 ^ n1270 ;
  assign n1091 = x29 ^ x13 ;
  assign n1092 = x157 ^ x141 ;
  assign n1264 = n1091 & n1092 ;
  assign n1089 = x28 ^ x12 ;
  assign n1090 = x156 ^ x140 ;
  assign n1263 = n1089 & n1090 ;
  assign n1268 = n1264 ^ n1263 ;
  assign n1289 = n1275 ^ n1268 ;
  assign n1087 = x27 ^ x11 ;
  assign n1088 = x155 ^ x139 ;
  assign n1239 = n1087 & n1088 ;
  assign n1085 = x26 ^ x10 ;
  assign n1086 = x154 ^ x138 ;
  assign n1238 = n1085 & n1086 ;
  assign n1243 = n1239 ^ n1238 ;
  assign n1083 = x25 ^ x9 ;
  assign n1084 = x153 ^ x137 ;
  assign n1232 = n1083 & n1084 ;
  assign n1081 = x24 ^ x8 ;
  assign n1082 = x152 ^ x136 ;
  assign n1231 = n1081 & n1082 ;
  assign n1236 = n1232 ^ n1231 ;
  assign n1257 = n1243 ^ n1236 ;
  assign n1338 = n1289 ^ n1257 ;
  assign n1079 = x23 ^ x7 ;
  assign n1080 = x151 ^ x135 ;
  assign n1152 = n1079 & n1080 ;
  assign n1077 = x22 ^ x6 ;
  assign n1078 = x150 ^ x134 ;
  assign n1151 = n1077 & n1078 ;
  assign n1156 = n1152 ^ n1151 ;
  assign n1075 = x21 ^ x5 ;
  assign n1076 = x149 ^ x133 ;
  assign n1145 = n1075 & n1076 ;
  assign n1073 = x20 ^ x4 ;
  assign n1074 = x148 ^ x132 ;
  assign n1144 = n1073 & n1074 ;
  assign n1149 = n1145 ^ n1144 ;
  assign n1170 = n1156 ^ n1149 ;
  assign n1071 = x19 ^ x3 ;
  assign n1072 = x147 ^ x131 ;
  assign n1120 = n1071 & n1072 ;
  assign n1069 = x18 ^ x2 ;
  assign n1070 = x146 ^ x130 ;
  assign n1119 = n1069 & n1070 ;
  assign n1124 = n1120 ^ n1119 ;
  assign n1067 = x17 ^ x1 ;
  assign n1068 = x145 ^ x129 ;
  assign n1113 = n1067 & n1068 ;
  assign n1065 = x16 ^ x0 ;
  assign n1066 = x144 ^ x128 ;
  assign n1112 = n1065 & n1066 ;
  assign n1117 = n1113 ^ n1112 ;
  assign n1138 = n1124 ^ n1117 ;
  assign n1219 = n1170 ^ n1138 ;
  assign n1492 = n1338 ^ n1219 ;
  assign n1532 = n1516 ^ n1492 ;
  assign n1533 = n1532 ^ n1050 ;
  assign n4289 = n2840 ^ n1533 ;
  assign n12800 = n8401 ^ n4289 ;
  assign n6691 = n6514 ^ n6512 ;
  assign n6692 = n6515 ^ n6513 ;
  assign n6693 = n6691 & n6692 ;
  assign n6695 = n6693 ^ n6689 ;
  assign n6684 = n6510 ^ n6508 ;
  assign n6685 = n6511 ^ n6509 ;
  assign n6686 = n6684 & n6685 ;
  assign n6688 = n6686 ^ n6682 ;
  assign n6709 = n6695 ^ n6688 ;
  assign n6659 = n6506 ^ n6504 ;
  assign n6660 = n6507 ^ n6505 ;
  assign n6661 = n6659 & n6660 ;
  assign n6663 = n6661 ^ n6657 ;
  assign n6652 = n6502 ^ n6500 ;
  assign n6653 = n6503 ^ n6501 ;
  assign n6654 = n6652 & n6653 ;
  assign n6656 = n6654 ^ n6650 ;
  assign n6677 = n6663 ^ n6656 ;
  assign n6758 = n6709 ^ n6677 ;
  assign n6572 = n6498 ^ n6496 ;
  assign n6573 = n6499 ^ n6497 ;
  assign n6574 = n6572 & n6573 ;
  assign n6576 = n6574 ^ n6570 ;
  assign n6565 = n6494 ^ n6492 ;
  assign n6566 = n6495 ^ n6493 ;
  assign n6567 = n6565 & n6566 ;
  assign n6569 = n6567 ^ n6563 ;
  assign n6590 = n6576 ^ n6569 ;
  assign n6540 = n6490 ^ n6488 ;
  assign n6541 = n6491 ^ n6489 ;
  assign n6542 = n6540 & n6541 ;
  assign n6544 = n6542 ^ n6538 ;
  assign n6533 = n6486 ^ n6484 ;
  assign n6534 = n6487 ^ n6485 ;
  assign n6535 = n6533 & n6534 ;
  assign n6537 = n6535 ^ n6531 ;
  assign n6558 = n6544 ^ n6537 ;
  assign n6639 = n6590 ^ n6558 ;
  assign n6912 = n6758 ^ n6639 ;
  assign n6953 = n6936 ^ n6912 ;
  assign n6954 = n6953 ^ n6471 ;
  assign n5384 = n5207 ^ n5205 ;
  assign n5385 = n5208 ^ n5206 ;
  assign n5386 = n5384 & n5385 ;
  assign n5388 = n5386 ^ n5382 ;
  assign n5377 = n5203 ^ n5201 ;
  assign n5378 = n5204 ^ n5202 ;
  assign n5379 = n5377 & n5378 ;
  assign n5381 = n5379 ^ n5375 ;
  assign n5402 = n5388 ^ n5381 ;
  assign n5352 = n5199 ^ n5197 ;
  assign n5353 = n5200 ^ n5198 ;
  assign n5354 = n5352 & n5353 ;
  assign n5356 = n5354 ^ n5350 ;
  assign n5345 = n5195 ^ n5193 ;
  assign n5346 = n5196 ^ n5194 ;
  assign n5347 = n5345 & n5346 ;
  assign n5349 = n5347 ^ n5343 ;
  assign n5370 = n5356 ^ n5349 ;
  assign n5451 = n5402 ^ n5370 ;
  assign n5265 = n5191 ^ n5189 ;
  assign n5266 = n5192 ^ n5190 ;
  assign n5267 = n5265 & n5266 ;
  assign n5269 = n5267 ^ n5263 ;
  assign n5258 = n5187 ^ n5185 ;
  assign n5259 = n5188 ^ n5186 ;
  assign n5260 = n5258 & n5259 ;
  assign n5262 = n5260 ^ n5256 ;
  assign n5283 = n5269 ^ n5262 ;
  assign n5233 = n5183 ^ n5181 ;
  assign n5234 = n5184 ^ n5182 ;
  assign n5235 = n5233 & n5234 ;
  assign n5237 = n5235 ^ n5231 ;
  assign n5226 = n5179 ^ n5177 ;
  assign n5227 = n5180 ^ n5178 ;
  assign n5228 = n5226 & n5227 ;
  assign n5230 = n5228 ^ n5224 ;
  assign n5251 = n5237 ^ n5230 ;
  assign n5332 = n5283 ^ n5251 ;
  assign n5605 = n5451 ^ n5332 ;
  assign n5646 = n5629 ^ n5605 ;
  assign n5647 = n5646 ^ n5164 ;
  assign n8402 = n6954 ^ n5647 ;
  assign n2579 = n2402 ^ n2400 ;
  assign n2580 = n2403 ^ n2401 ;
  assign n2581 = n2579 & n2580 ;
  assign n2583 = n2581 ^ n2577 ;
  assign n2572 = n2398 ^ n2396 ;
  assign n2573 = n2399 ^ n2397 ;
  assign n2574 = n2572 & n2573 ;
  assign n2576 = n2574 ^ n2570 ;
  assign n2597 = n2583 ^ n2576 ;
  assign n2547 = n2394 ^ n2392 ;
  assign n2548 = n2395 ^ n2393 ;
  assign n2549 = n2547 & n2548 ;
  assign n2551 = n2549 ^ n2545 ;
  assign n2540 = n2390 ^ n2388 ;
  assign n2541 = n2391 ^ n2389 ;
  assign n2542 = n2540 & n2541 ;
  assign n2544 = n2542 ^ n2538 ;
  assign n2565 = n2551 ^ n2544 ;
  assign n2646 = n2597 ^ n2565 ;
  assign n2460 = n2386 ^ n2384 ;
  assign n2461 = n2387 ^ n2385 ;
  assign n2462 = n2460 & n2461 ;
  assign n2464 = n2462 ^ n2458 ;
  assign n2453 = n2382 ^ n2380 ;
  assign n2454 = n2383 ^ n2381 ;
  assign n2455 = n2453 & n2454 ;
  assign n2457 = n2455 ^ n2451 ;
  assign n2478 = n2464 ^ n2457 ;
  assign n2428 = n2378 ^ n2376 ;
  assign n2429 = n2379 ^ n2377 ;
  assign n2430 = n2428 & n2429 ;
  assign n2432 = n2430 ^ n2426 ;
  assign n2421 = n2374 ^ n2372 ;
  assign n2422 = n2375 ^ n2373 ;
  assign n2423 = n2421 & n2422 ;
  assign n2425 = n2423 ^ n2419 ;
  assign n2446 = n2432 ^ n2425 ;
  assign n2527 = n2478 ^ n2446 ;
  assign n2800 = n2646 ^ n2527 ;
  assign n2841 = n2824 ^ n2800 ;
  assign n2842 = n2841 ^ n2359 ;
  assign n1272 = n1095 ^ n1093 ;
  assign n1273 = n1096 ^ n1094 ;
  assign n1274 = n1272 & n1273 ;
  assign n1276 = n1274 ^ n1270 ;
  assign n1265 = n1091 ^ n1089 ;
  assign n1266 = n1092 ^ n1090 ;
  assign n1267 = n1265 & n1266 ;
  assign n1269 = n1267 ^ n1263 ;
  assign n1290 = n1276 ^ n1269 ;
  assign n1240 = n1087 ^ n1085 ;
  assign n1241 = n1088 ^ n1086 ;
  assign n1242 = n1240 & n1241 ;
  assign n1244 = n1242 ^ n1238 ;
  assign n1233 = n1083 ^ n1081 ;
  assign n1234 = n1084 ^ n1082 ;
  assign n1235 = n1233 & n1234 ;
  assign n1237 = n1235 ^ n1231 ;
  assign n1258 = n1244 ^ n1237 ;
  assign n1339 = n1290 ^ n1258 ;
  assign n1153 = n1079 ^ n1077 ;
  assign n1154 = n1080 ^ n1078 ;
  assign n1155 = n1153 & n1154 ;
  assign n1157 = n1155 ^ n1151 ;
  assign n1146 = n1075 ^ n1073 ;
  assign n1147 = n1076 ^ n1074 ;
  assign n1148 = n1146 & n1147 ;
  assign n1150 = n1148 ^ n1144 ;
  assign n1171 = n1157 ^ n1150 ;
  assign n1121 = n1071 ^ n1069 ;
  assign n1122 = n1072 ^ n1070 ;
  assign n1123 = n1121 & n1122 ;
  assign n1125 = n1123 ^ n1119 ;
  assign n1114 = n1067 ^ n1065 ;
  assign n1115 = n1068 ^ n1066 ;
  assign n1116 = n1114 & n1115 ;
  assign n1118 = n1116 ^ n1112 ;
  assign n1139 = n1125 ^ n1118 ;
  assign n1220 = n1171 ^ n1139 ;
  assign n1493 = n1339 ^ n1220 ;
  assign n1534 = n1517 ^ n1493 ;
  assign n1535 = n1534 ^ n1052 ;
  assign n4290 = n2842 ^ n1535 ;
  assign n12801 = n8402 ^ n4290 ;
  assign n6698 = n6514 ^ n6510 ;
  assign n6699 = n6515 ^ n6511 ;
  assign n6702 = n6698 & n6699 ;
  assign n6696 = n6512 ^ n6508 ;
  assign n6697 = n6513 ^ n6509 ;
  assign n6701 = n6696 & n6697 ;
  assign n6706 = n6702 ^ n6701 ;
  assign n6710 = n6708 ^ n6706 ;
  assign n6711 = n6710 ^ n6695 ;
  assign n6666 = n6506 ^ n6502 ;
  assign n6667 = n6507 ^ n6503 ;
  assign n6670 = n6666 & n6667 ;
  assign n6664 = n6504 ^ n6500 ;
  assign n6665 = n6505 ^ n6501 ;
  assign n6669 = n6664 & n6665 ;
  assign n6674 = n6670 ^ n6669 ;
  assign n6678 = n6676 ^ n6674 ;
  assign n6679 = n6678 ^ n6663 ;
  assign n6759 = n6711 ^ n6679 ;
  assign n6579 = n6498 ^ n6494 ;
  assign n6580 = n6499 ^ n6495 ;
  assign n6583 = n6579 & n6580 ;
  assign n6577 = n6496 ^ n6492 ;
  assign n6578 = n6497 ^ n6493 ;
  assign n6582 = n6577 & n6578 ;
  assign n6587 = n6583 ^ n6582 ;
  assign n6591 = n6589 ^ n6587 ;
  assign n6592 = n6591 ^ n6576 ;
  assign n6547 = n6490 ^ n6486 ;
  assign n6548 = n6491 ^ n6487 ;
  assign n6551 = n6547 & n6548 ;
  assign n6545 = n6488 ^ n6484 ;
  assign n6546 = n6489 ^ n6485 ;
  assign n6550 = n6545 & n6546 ;
  assign n6555 = n6551 ^ n6550 ;
  assign n6559 = n6557 ^ n6555 ;
  assign n6560 = n6559 ^ n6544 ;
  assign n6640 = n6592 ^ n6560 ;
  assign n6913 = n6759 ^ n6640 ;
  assign n6955 = n6937 ^ n6913 ;
  assign n6956 = n6955 ^ n6473 ;
  assign n5391 = n5207 ^ n5203 ;
  assign n5392 = n5208 ^ n5204 ;
  assign n5395 = n5391 & n5392 ;
  assign n5389 = n5205 ^ n5201 ;
  assign n5390 = n5206 ^ n5202 ;
  assign n5394 = n5389 & n5390 ;
  assign n5399 = n5395 ^ n5394 ;
  assign n5403 = n5401 ^ n5399 ;
  assign n5404 = n5403 ^ n5388 ;
  assign n5359 = n5199 ^ n5195 ;
  assign n5360 = n5200 ^ n5196 ;
  assign n5363 = n5359 & n5360 ;
  assign n5357 = n5197 ^ n5193 ;
  assign n5358 = n5198 ^ n5194 ;
  assign n5362 = n5357 & n5358 ;
  assign n5367 = n5363 ^ n5362 ;
  assign n5371 = n5369 ^ n5367 ;
  assign n5372 = n5371 ^ n5356 ;
  assign n5452 = n5404 ^ n5372 ;
  assign n5272 = n5191 ^ n5187 ;
  assign n5273 = n5192 ^ n5188 ;
  assign n5276 = n5272 & n5273 ;
  assign n5270 = n5189 ^ n5185 ;
  assign n5271 = n5190 ^ n5186 ;
  assign n5275 = n5270 & n5271 ;
  assign n5280 = n5276 ^ n5275 ;
  assign n5284 = n5282 ^ n5280 ;
  assign n5285 = n5284 ^ n5269 ;
  assign n5240 = n5183 ^ n5179 ;
  assign n5241 = n5184 ^ n5180 ;
  assign n5244 = n5240 & n5241 ;
  assign n5238 = n5181 ^ n5177 ;
  assign n5239 = n5182 ^ n5178 ;
  assign n5243 = n5238 & n5239 ;
  assign n5248 = n5244 ^ n5243 ;
  assign n5252 = n5250 ^ n5248 ;
  assign n5253 = n5252 ^ n5237 ;
  assign n5333 = n5285 ^ n5253 ;
  assign n5606 = n5452 ^ n5333 ;
  assign n5648 = n5630 ^ n5606 ;
  assign n5649 = n5648 ^ n5166 ;
  assign n8403 = n6956 ^ n5649 ;
  assign n2586 = n2402 ^ n2398 ;
  assign n2587 = n2403 ^ n2399 ;
  assign n2590 = n2586 & n2587 ;
  assign n2584 = n2400 ^ n2396 ;
  assign n2585 = n2401 ^ n2397 ;
  assign n2589 = n2584 & n2585 ;
  assign n2594 = n2590 ^ n2589 ;
  assign n2598 = n2596 ^ n2594 ;
  assign n2599 = n2598 ^ n2583 ;
  assign n2554 = n2394 ^ n2390 ;
  assign n2555 = n2395 ^ n2391 ;
  assign n2558 = n2554 & n2555 ;
  assign n2552 = n2392 ^ n2388 ;
  assign n2553 = n2393 ^ n2389 ;
  assign n2557 = n2552 & n2553 ;
  assign n2562 = n2558 ^ n2557 ;
  assign n2566 = n2564 ^ n2562 ;
  assign n2567 = n2566 ^ n2551 ;
  assign n2647 = n2599 ^ n2567 ;
  assign n2467 = n2386 ^ n2382 ;
  assign n2468 = n2387 ^ n2383 ;
  assign n2471 = n2467 & n2468 ;
  assign n2465 = n2384 ^ n2380 ;
  assign n2466 = n2385 ^ n2381 ;
  assign n2470 = n2465 & n2466 ;
  assign n2475 = n2471 ^ n2470 ;
  assign n2479 = n2477 ^ n2475 ;
  assign n2480 = n2479 ^ n2464 ;
  assign n2435 = n2378 ^ n2374 ;
  assign n2436 = n2379 ^ n2375 ;
  assign n2439 = n2435 & n2436 ;
  assign n2433 = n2376 ^ n2372 ;
  assign n2434 = n2377 ^ n2373 ;
  assign n2438 = n2433 & n2434 ;
  assign n2443 = n2439 ^ n2438 ;
  assign n2447 = n2445 ^ n2443 ;
  assign n2448 = n2447 ^ n2432 ;
  assign n2528 = n2480 ^ n2448 ;
  assign n2801 = n2647 ^ n2528 ;
  assign n2843 = n2825 ^ n2801 ;
  assign n2844 = n2843 ^ n2361 ;
  assign n1279 = n1095 ^ n1091 ;
  assign n1280 = n1096 ^ n1092 ;
  assign n1283 = n1279 & n1280 ;
  assign n1277 = n1093 ^ n1089 ;
  assign n1278 = n1094 ^ n1090 ;
  assign n1282 = n1277 & n1278 ;
  assign n1287 = n1283 ^ n1282 ;
  assign n1291 = n1289 ^ n1287 ;
  assign n1292 = n1291 ^ n1276 ;
  assign n1247 = n1087 ^ n1083 ;
  assign n1248 = n1088 ^ n1084 ;
  assign n1251 = n1247 & n1248 ;
  assign n1245 = n1085 ^ n1081 ;
  assign n1246 = n1086 ^ n1082 ;
  assign n1250 = n1245 & n1246 ;
  assign n1255 = n1251 ^ n1250 ;
  assign n1259 = n1257 ^ n1255 ;
  assign n1260 = n1259 ^ n1244 ;
  assign n1340 = n1292 ^ n1260 ;
  assign n1160 = n1079 ^ n1075 ;
  assign n1161 = n1080 ^ n1076 ;
  assign n1164 = n1160 & n1161 ;
  assign n1158 = n1077 ^ n1073 ;
  assign n1159 = n1078 ^ n1074 ;
  assign n1163 = n1158 & n1159 ;
  assign n1168 = n1164 ^ n1163 ;
  assign n1172 = n1170 ^ n1168 ;
  assign n1173 = n1172 ^ n1157 ;
  assign n1128 = n1071 ^ n1067 ;
  assign n1129 = n1072 ^ n1068 ;
  assign n1132 = n1128 & n1129 ;
  assign n1126 = n1069 ^ n1065 ;
  assign n1127 = n1070 ^ n1066 ;
  assign n1131 = n1126 & n1127 ;
  assign n1136 = n1132 ^ n1131 ;
  assign n1140 = n1138 ^ n1136 ;
  assign n1141 = n1140 ^ n1125 ;
  assign n1221 = n1173 ^ n1141 ;
  assign n1494 = n1340 ^ n1221 ;
  assign n1536 = n1518 ^ n1494 ;
  assign n1537 = n1536 ^ n1054 ;
  assign n4291 = n2844 ^ n1537 ;
  assign n12802 = n8403 ^ n4291 ;
  assign n6703 = n6698 ^ n6696 ;
  assign n6704 = n6699 ^ n6697 ;
  assign n6705 = n6703 & n6704 ;
  assign n6707 = n6705 ^ n6701 ;
  assign n6712 = n6709 ^ n6707 ;
  assign n6700 = n6695 ^ n6694 ;
  assign n6713 = n6712 ^ n6700 ;
  assign n6671 = n6666 ^ n6664 ;
  assign n6672 = n6667 ^ n6665 ;
  assign n6673 = n6671 & n6672 ;
  assign n6675 = n6673 ^ n6669 ;
  assign n6680 = n6677 ^ n6675 ;
  assign n6668 = n6663 ^ n6662 ;
  assign n6681 = n6680 ^ n6668 ;
  assign n6760 = n6713 ^ n6681 ;
  assign n6584 = n6579 ^ n6577 ;
  assign n6585 = n6580 ^ n6578 ;
  assign n6586 = n6584 & n6585 ;
  assign n6588 = n6586 ^ n6582 ;
  assign n6593 = n6590 ^ n6588 ;
  assign n6581 = n6576 ^ n6575 ;
  assign n6594 = n6593 ^ n6581 ;
  assign n6552 = n6547 ^ n6545 ;
  assign n6553 = n6548 ^ n6546 ;
  assign n6554 = n6552 & n6553 ;
  assign n6556 = n6554 ^ n6550 ;
  assign n6561 = n6558 ^ n6556 ;
  assign n6549 = n6544 ^ n6543 ;
  assign n6562 = n6561 ^ n6549 ;
  assign n6641 = n6594 ^ n6562 ;
  assign n6914 = n6760 ^ n6641 ;
  assign n6957 = n6938 ^ n6914 ;
  assign n6958 = n6957 ^ n6475 ;
  assign n5396 = n5391 ^ n5389 ;
  assign n5397 = n5392 ^ n5390 ;
  assign n5398 = n5396 & n5397 ;
  assign n5400 = n5398 ^ n5394 ;
  assign n5405 = n5402 ^ n5400 ;
  assign n5393 = n5388 ^ n5387 ;
  assign n5406 = n5405 ^ n5393 ;
  assign n5364 = n5359 ^ n5357 ;
  assign n5365 = n5360 ^ n5358 ;
  assign n5366 = n5364 & n5365 ;
  assign n5368 = n5366 ^ n5362 ;
  assign n5373 = n5370 ^ n5368 ;
  assign n5361 = n5356 ^ n5355 ;
  assign n5374 = n5373 ^ n5361 ;
  assign n5453 = n5406 ^ n5374 ;
  assign n5277 = n5272 ^ n5270 ;
  assign n5278 = n5273 ^ n5271 ;
  assign n5279 = n5277 & n5278 ;
  assign n5281 = n5279 ^ n5275 ;
  assign n5286 = n5283 ^ n5281 ;
  assign n5274 = n5269 ^ n5268 ;
  assign n5287 = n5286 ^ n5274 ;
  assign n5245 = n5240 ^ n5238 ;
  assign n5246 = n5241 ^ n5239 ;
  assign n5247 = n5245 & n5246 ;
  assign n5249 = n5247 ^ n5243 ;
  assign n5254 = n5251 ^ n5249 ;
  assign n5242 = n5237 ^ n5236 ;
  assign n5255 = n5254 ^ n5242 ;
  assign n5334 = n5287 ^ n5255 ;
  assign n5607 = n5453 ^ n5334 ;
  assign n5650 = n5631 ^ n5607 ;
  assign n5651 = n5650 ^ n5168 ;
  assign n8404 = n6958 ^ n5651 ;
  assign n2591 = n2586 ^ n2584 ;
  assign n2592 = n2587 ^ n2585 ;
  assign n2593 = n2591 & n2592 ;
  assign n2595 = n2593 ^ n2589 ;
  assign n2600 = n2597 ^ n2595 ;
  assign n2588 = n2583 ^ n2582 ;
  assign n2601 = n2600 ^ n2588 ;
  assign n2559 = n2554 ^ n2552 ;
  assign n2560 = n2555 ^ n2553 ;
  assign n2561 = n2559 & n2560 ;
  assign n2563 = n2561 ^ n2557 ;
  assign n2568 = n2565 ^ n2563 ;
  assign n2556 = n2551 ^ n2550 ;
  assign n2569 = n2568 ^ n2556 ;
  assign n2648 = n2601 ^ n2569 ;
  assign n2472 = n2467 ^ n2465 ;
  assign n2473 = n2468 ^ n2466 ;
  assign n2474 = n2472 & n2473 ;
  assign n2476 = n2474 ^ n2470 ;
  assign n2481 = n2478 ^ n2476 ;
  assign n2469 = n2464 ^ n2463 ;
  assign n2482 = n2481 ^ n2469 ;
  assign n2440 = n2435 ^ n2433 ;
  assign n2441 = n2436 ^ n2434 ;
  assign n2442 = n2440 & n2441 ;
  assign n2444 = n2442 ^ n2438 ;
  assign n2449 = n2446 ^ n2444 ;
  assign n2437 = n2432 ^ n2431 ;
  assign n2450 = n2449 ^ n2437 ;
  assign n2529 = n2482 ^ n2450 ;
  assign n2802 = n2648 ^ n2529 ;
  assign n2845 = n2826 ^ n2802 ;
  assign n2846 = n2845 ^ n2363 ;
  assign n1284 = n1279 ^ n1277 ;
  assign n1285 = n1280 ^ n1278 ;
  assign n1286 = n1284 & n1285 ;
  assign n1288 = n1286 ^ n1282 ;
  assign n1293 = n1290 ^ n1288 ;
  assign n1281 = n1276 ^ n1275 ;
  assign n1294 = n1293 ^ n1281 ;
  assign n1252 = n1247 ^ n1245 ;
  assign n1253 = n1248 ^ n1246 ;
  assign n1254 = n1252 & n1253 ;
  assign n1256 = n1254 ^ n1250 ;
  assign n1261 = n1258 ^ n1256 ;
  assign n1249 = n1244 ^ n1243 ;
  assign n1262 = n1261 ^ n1249 ;
  assign n1341 = n1294 ^ n1262 ;
  assign n1165 = n1160 ^ n1158 ;
  assign n1166 = n1161 ^ n1159 ;
  assign n1167 = n1165 & n1166 ;
  assign n1169 = n1167 ^ n1163 ;
  assign n1174 = n1171 ^ n1169 ;
  assign n1162 = n1157 ^ n1156 ;
  assign n1175 = n1174 ^ n1162 ;
  assign n1133 = n1128 ^ n1126 ;
  assign n1134 = n1129 ^ n1127 ;
  assign n1135 = n1133 & n1134 ;
  assign n1137 = n1135 ^ n1131 ;
  assign n1142 = n1139 ^ n1137 ;
  assign n1130 = n1125 ^ n1124 ;
  assign n1143 = n1142 ^ n1130 ;
  assign n1222 = n1175 ^ n1143 ;
  assign n1495 = n1341 ^ n1222 ;
  assign n1538 = n1519 ^ n1495 ;
  assign n1539 = n1538 ^ n1056 ;
  assign n4292 = n2846 ^ n1539 ;
  assign n12803 = n8404 ^ n4292 ;
  assign n6720 = n6514 ^ n6506 ;
  assign n6721 = n6515 ^ n6507 ;
  assign n6733 = n6720 & n6721 ;
  assign n6718 = n6512 ^ n6504 ;
  assign n6719 = n6513 ^ n6505 ;
  assign n6732 = n6718 & n6719 ;
  assign n6737 = n6733 ^ n6732 ;
  assign n6716 = n6510 ^ n6502 ;
  assign n6717 = n6511 ^ n6503 ;
  assign n6726 = n6716 & n6717 ;
  assign n6714 = n6508 ^ n6500 ;
  assign n6715 = n6509 ^ n6501 ;
  assign n6725 = n6714 & n6715 ;
  assign n6730 = n6726 ^ n6725 ;
  assign n6751 = n6737 ^ n6730 ;
  assign n6761 = n6757 ^ n6751 ;
  assign n6762 = n6761 ^ n6711 ;
  assign n6601 = n6498 ^ n6490 ;
  assign n6602 = n6499 ^ n6491 ;
  assign n6614 = n6601 & n6602 ;
  assign n6599 = n6496 ^ n6488 ;
  assign n6600 = n6497 ^ n6489 ;
  assign n6613 = n6599 & n6600 ;
  assign n6618 = n6614 ^ n6613 ;
  assign n6597 = n6494 ^ n6486 ;
  assign n6598 = n6495 ^ n6487 ;
  assign n6607 = n6597 & n6598 ;
  assign n6595 = n6492 ^ n6484 ;
  assign n6596 = n6493 ^ n6485 ;
  assign n6606 = n6595 & n6596 ;
  assign n6611 = n6607 ^ n6606 ;
  assign n6632 = n6618 ^ n6611 ;
  assign n6642 = n6638 ^ n6632 ;
  assign n6643 = n6642 ^ n6592 ;
  assign n6915 = n6762 ^ n6643 ;
  assign n6959 = n6939 ^ n6915 ;
  assign n6960 = n6959 ^ n6477 ;
  assign n5413 = n5207 ^ n5199 ;
  assign n5414 = n5208 ^ n5200 ;
  assign n5426 = n5413 & n5414 ;
  assign n5411 = n5205 ^ n5197 ;
  assign n5412 = n5206 ^ n5198 ;
  assign n5425 = n5411 & n5412 ;
  assign n5430 = n5426 ^ n5425 ;
  assign n5409 = n5203 ^ n5195 ;
  assign n5410 = n5204 ^ n5196 ;
  assign n5419 = n5409 & n5410 ;
  assign n5407 = n5201 ^ n5193 ;
  assign n5408 = n5202 ^ n5194 ;
  assign n5418 = n5407 & n5408 ;
  assign n5423 = n5419 ^ n5418 ;
  assign n5444 = n5430 ^ n5423 ;
  assign n5454 = n5450 ^ n5444 ;
  assign n5455 = n5454 ^ n5404 ;
  assign n5294 = n5191 ^ n5183 ;
  assign n5295 = n5192 ^ n5184 ;
  assign n5307 = n5294 & n5295 ;
  assign n5292 = n5189 ^ n5181 ;
  assign n5293 = n5190 ^ n5182 ;
  assign n5306 = n5292 & n5293 ;
  assign n5311 = n5307 ^ n5306 ;
  assign n5290 = n5187 ^ n5179 ;
  assign n5291 = n5188 ^ n5180 ;
  assign n5300 = n5290 & n5291 ;
  assign n5288 = n5185 ^ n5177 ;
  assign n5289 = n5186 ^ n5178 ;
  assign n5299 = n5288 & n5289 ;
  assign n5304 = n5300 ^ n5299 ;
  assign n5325 = n5311 ^ n5304 ;
  assign n5335 = n5331 ^ n5325 ;
  assign n5336 = n5335 ^ n5285 ;
  assign n5608 = n5455 ^ n5336 ;
  assign n5652 = n5632 ^ n5608 ;
  assign n5653 = n5652 ^ n5170 ;
  assign n8405 = n6960 ^ n5653 ;
  assign n2608 = n2402 ^ n2394 ;
  assign n2609 = n2403 ^ n2395 ;
  assign n2621 = n2608 & n2609 ;
  assign n2606 = n2400 ^ n2392 ;
  assign n2607 = n2401 ^ n2393 ;
  assign n2620 = n2606 & n2607 ;
  assign n2625 = n2621 ^ n2620 ;
  assign n2604 = n2398 ^ n2390 ;
  assign n2605 = n2399 ^ n2391 ;
  assign n2614 = n2604 & n2605 ;
  assign n2602 = n2396 ^ n2388 ;
  assign n2603 = n2397 ^ n2389 ;
  assign n2613 = n2602 & n2603 ;
  assign n2618 = n2614 ^ n2613 ;
  assign n2639 = n2625 ^ n2618 ;
  assign n2649 = n2645 ^ n2639 ;
  assign n2650 = n2649 ^ n2599 ;
  assign n2489 = n2386 ^ n2378 ;
  assign n2490 = n2387 ^ n2379 ;
  assign n2502 = n2489 & n2490 ;
  assign n2487 = n2384 ^ n2376 ;
  assign n2488 = n2385 ^ n2377 ;
  assign n2501 = n2487 & n2488 ;
  assign n2506 = n2502 ^ n2501 ;
  assign n2485 = n2382 ^ n2374 ;
  assign n2486 = n2383 ^ n2375 ;
  assign n2495 = n2485 & n2486 ;
  assign n2483 = n2380 ^ n2372 ;
  assign n2484 = n2381 ^ n2373 ;
  assign n2494 = n2483 & n2484 ;
  assign n2499 = n2495 ^ n2494 ;
  assign n2520 = n2506 ^ n2499 ;
  assign n2530 = n2526 ^ n2520 ;
  assign n2531 = n2530 ^ n2480 ;
  assign n2803 = n2650 ^ n2531 ;
  assign n2847 = n2827 ^ n2803 ;
  assign n2848 = n2847 ^ n2365 ;
  assign n1301 = n1095 ^ n1087 ;
  assign n1302 = n1096 ^ n1088 ;
  assign n1314 = n1301 & n1302 ;
  assign n1299 = n1093 ^ n1085 ;
  assign n1300 = n1094 ^ n1086 ;
  assign n1313 = n1299 & n1300 ;
  assign n1318 = n1314 ^ n1313 ;
  assign n1297 = n1091 ^ n1083 ;
  assign n1298 = n1092 ^ n1084 ;
  assign n1307 = n1297 & n1298 ;
  assign n1295 = n1089 ^ n1081 ;
  assign n1296 = n1090 ^ n1082 ;
  assign n1306 = n1295 & n1296 ;
  assign n1311 = n1307 ^ n1306 ;
  assign n1332 = n1318 ^ n1311 ;
  assign n1342 = n1338 ^ n1332 ;
  assign n1343 = n1342 ^ n1292 ;
  assign n1182 = n1079 ^ n1071 ;
  assign n1183 = n1080 ^ n1072 ;
  assign n1195 = n1182 & n1183 ;
  assign n1180 = n1077 ^ n1069 ;
  assign n1181 = n1078 ^ n1070 ;
  assign n1194 = n1180 & n1181 ;
  assign n1199 = n1195 ^ n1194 ;
  assign n1178 = n1075 ^ n1067 ;
  assign n1179 = n1076 ^ n1068 ;
  assign n1188 = n1178 & n1179 ;
  assign n1176 = n1073 ^ n1065 ;
  assign n1177 = n1074 ^ n1066 ;
  assign n1187 = n1176 & n1177 ;
  assign n1192 = n1188 ^ n1187 ;
  assign n1213 = n1199 ^ n1192 ;
  assign n1223 = n1219 ^ n1213 ;
  assign n1224 = n1223 ^ n1173 ;
  assign n1496 = n1343 ^ n1224 ;
  assign n1540 = n1520 ^ n1496 ;
  assign n1541 = n1540 ^ n1058 ;
  assign n4293 = n2848 ^ n1541 ;
  assign n12804 = n8405 ^ n4293 ;
  assign n6734 = n6720 ^ n6718 ;
  assign n6735 = n6721 ^ n6719 ;
  assign n6736 = n6734 & n6735 ;
  assign n6738 = n6736 ^ n6732 ;
  assign n6727 = n6716 ^ n6714 ;
  assign n6728 = n6717 ^ n6715 ;
  assign n6729 = n6727 & n6728 ;
  assign n6731 = n6729 ^ n6725 ;
  assign n6752 = n6738 ^ n6731 ;
  assign n6763 = n6758 ^ n6752 ;
  assign n6764 = n6763 ^ n6713 ;
  assign n6615 = n6601 ^ n6599 ;
  assign n6616 = n6602 ^ n6600 ;
  assign n6617 = n6615 & n6616 ;
  assign n6619 = n6617 ^ n6613 ;
  assign n6608 = n6597 ^ n6595 ;
  assign n6609 = n6598 ^ n6596 ;
  assign n6610 = n6608 & n6609 ;
  assign n6612 = n6610 ^ n6606 ;
  assign n6633 = n6619 ^ n6612 ;
  assign n6644 = n6639 ^ n6633 ;
  assign n6645 = n6644 ^ n6594 ;
  assign n6916 = n6764 ^ n6645 ;
  assign n6961 = n6940 ^ n6916 ;
  assign n6962 = n6961 ^ n6479 ;
  assign n5427 = n5413 ^ n5411 ;
  assign n5428 = n5414 ^ n5412 ;
  assign n5429 = n5427 & n5428 ;
  assign n5431 = n5429 ^ n5425 ;
  assign n5420 = n5409 ^ n5407 ;
  assign n5421 = n5410 ^ n5408 ;
  assign n5422 = n5420 & n5421 ;
  assign n5424 = n5422 ^ n5418 ;
  assign n5445 = n5431 ^ n5424 ;
  assign n5456 = n5451 ^ n5445 ;
  assign n5457 = n5456 ^ n5406 ;
  assign n5308 = n5294 ^ n5292 ;
  assign n5309 = n5295 ^ n5293 ;
  assign n5310 = n5308 & n5309 ;
  assign n5312 = n5310 ^ n5306 ;
  assign n5301 = n5290 ^ n5288 ;
  assign n5302 = n5291 ^ n5289 ;
  assign n5303 = n5301 & n5302 ;
  assign n5305 = n5303 ^ n5299 ;
  assign n5326 = n5312 ^ n5305 ;
  assign n5337 = n5332 ^ n5326 ;
  assign n5338 = n5337 ^ n5287 ;
  assign n5609 = n5457 ^ n5338 ;
  assign n5654 = n5633 ^ n5609 ;
  assign n5655 = n5654 ^ n5172 ;
  assign n8406 = n6962 ^ n5655 ;
  assign n2622 = n2608 ^ n2606 ;
  assign n2623 = n2609 ^ n2607 ;
  assign n2624 = n2622 & n2623 ;
  assign n2626 = n2624 ^ n2620 ;
  assign n2615 = n2604 ^ n2602 ;
  assign n2616 = n2605 ^ n2603 ;
  assign n2617 = n2615 & n2616 ;
  assign n2619 = n2617 ^ n2613 ;
  assign n2640 = n2626 ^ n2619 ;
  assign n2651 = n2646 ^ n2640 ;
  assign n2652 = n2651 ^ n2601 ;
  assign n2503 = n2489 ^ n2487 ;
  assign n2504 = n2490 ^ n2488 ;
  assign n2505 = n2503 & n2504 ;
  assign n2507 = n2505 ^ n2501 ;
  assign n2496 = n2485 ^ n2483 ;
  assign n2497 = n2486 ^ n2484 ;
  assign n2498 = n2496 & n2497 ;
  assign n2500 = n2498 ^ n2494 ;
  assign n2521 = n2507 ^ n2500 ;
  assign n2532 = n2527 ^ n2521 ;
  assign n2533 = n2532 ^ n2482 ;
  assign n2804 = n2652 ^ n2533 ;
  assign n2849 = n2828 ^ n2804 ;
  assign n2850 = n2849 ^ n2367 ;
  assign n1315 = n1301 ^ n1299 ;
  assign n1316 = n1302 ^ n1300 ;
  assign n1317 = n1315 & n1316 ;
  assign n1319 = n1317 ^ n1313 ;
  assign n1308 = n1297 ^ n1295 ;
  assign n1309 = n1298 ^ n1296 ;
  assign n1310 = n1308 & n1309 ;
  assign n1312 = n1310 ^ n1306 ;
  assign n1333 = n1319 ^ n1312 ;
  assign n1344 = n1339 ^ n1333 ;
  assign n1345 = n1344 ^ n1294 ;
  assign n1196 = n1182 ^ n1180 ;
  assign n1197 = n1183 ^ n1181 ;
  assign n1198 = n1196 & n1197 ;
  assign n1200 = n1198 ^ n1194 ;
  assign n1189 = n1178 ^ n1176 ;
  assign n1190 = n1179 ^ n1177 ;
  assign n1191 = n1189 & n1190 ;
  assign n1193 = n1191 ^ n1187 ;
  assign n1214 = n1200 ^ n1193 ;
  assign n1225 = n1220 ^ n1214 ;
  assign n1226 = n1225 ^ n1175 ;
  assign n1497 = n1345 ^ n1226 ;
  assign n1542 = n1521 ^ n1497 ;
  assign n1543 = n1542 ^ n1060 ;
  assign n4294 = n2850 ^ n1543 ;
  assign n12805 = n8406 ^ n4294 ;
  assign n6741 = n6720 ^ n6716 ;
  assign n6742 = n6721 ^ n6717 ;
  assign n6745 = n6741 & n6742 ;
  assign n6739 = n6718 ^ n6714 ;
  assign n6740 = n6719 ^ n6715 ;
  assign n6744 = n6739 & n6740 ;
  assign n6749 = n6745 ^ n6744 ;
  assign n6753 = n6751 ^ n6749 ;
  assign n6754 = n6753 ^ n6738 ;
  assign n6765 = n6759 ^ n6754 ;
  assign n6723 = n6713 ^ n6708 ;
  assign n6766 = n6765 ^ n6723 ;
  assign n6622 = n6601 ^ n6597 ;
  assign n6623 = n6602 ^ n6598 ;
  assign n6626 = n6622 & n6623 ;
  assign n6620 = n6599 ^ n6595 ;
  assign n6621 = n6600 ^ n6596 ;
  assign n6625 = n6620 & n6621 ;
  assign n6630 = n6626 ^ n6625 ;
  assign n6634 = n6632 ^ n6630 ;
  assign n6635 = n6634 ^ n6619 ;
  assign n6646 = n6640 ^ n6635 ;
  assign n6604 = n6594 ^ n6589 ;
  assign n6647 = n6646 ^ n6604 ;
  assign n6917 = n6766 ^ n6647 ;
  assign n6963 = n6941 ^ n6917 ;
  assign n6964 = n6963 ^ n6481 ;
  assign n5434 = n5413 ^ n5409 ;
  assign n5435 = n5414 ^ n5410 ;
  assign n5438 = n5434 & n5435 ;
  assign n5432 = n5411 ^ n5407 ;
  assign n5433 = n5412 ^ n5408 ;
  assign n5437 = n5432 & n5433 ;
  assign n5442 = n5438 ^ n5437 ;
  assign n5446 = n5444 ^ n5442 ;
  assign n5447 = n5446 ^ n5431 ;
  assign n5458 = n5452 ^ n5447 ;
  assign n5416 = n5406 ^ n5401 ;
  assign n5459 = n5458 ^ n5416 ;
  assign n5315 = n5294 ^ n5290 ;
  assign n5316 = n5295 ^ n5291 ;
  assign n5319 = n5315 & n5316 ;
  assign n5313 = n5292 ^ n5288 ;
  assign n5314 = n5293 ^ n5289 ;
  assign n5318 = n5313 & n5314 ;
  assign n5323 = n5319 ^ n5318 ;
  assign n5327 = n5325 ^ n5323 ;
  assign n5328 = n5327 ^ n5312 ;
  assign n5339 = n5333 ^ n5328 ;
  assign n5297 = n5287 ^ n5282 ;
  assign n5340 = n5339 ^ n5297 ;
  assign n5610 = n5459 ^ n5340 ;
  assign n5656 = n5634 ^ n5610 ;
  assign n5657 = n5656 ^ n5174 ;
  assign n8407 = n6964 ^ n5657 ;
  assign n2629 = n2608 ^ n2604 ;
  assign n2630 = n2609 ^ n2605 ;
  assign n2633 = n2629 & n2630 ;
  assign n2627 = n2606 ^ n2602 ;
  assign n2628 = n2607 ^ n2603 ;
  assign n2632 = n2627 & n2628 ;
  assign n2637 = n2633 ^ n2632 ;
  assign n2641 = n2639 ^ n2637 ;
  assign n2642 = n2641 ^ n2626 ;
  assign n2653 = n2647 ^ n2642 ;
  assign n2611 = n2601 ^ n2596 ;
  assign n2654 = n2653 ^ n2611 ;
  assign n2510 = n2489 ^ n2485 ;
  assign n2511 = n2490 ^ n2486 ;
  assign n2514 = n2510 & n2511 ;
  assign n2508 = n2487 ^ n2483 ;
  assign n2509 = n2488 ^ n2484 ;
  assign n2513 = n2508 & n2509 ;
  assign n2518 = n2514 ^ n2513 ;
  assign n2522 = n2520 ^ n2518 ;
  assign n2523 = n2522 ^ n2507 ;
  assign n2534 = n2528 ^ n2523 ;
  assign n2492 = n2482 ^ n2477 ;
  assign n2535 = n2534 ^ n2492 ;
  assign n2805 = n2654 ^ n2535 ;
  assign n2851 = n2829 ^ n2805 ;
  assign n2852 = n2851 ^ n2369 ;
  assign n1322 = n1301 ^ n1297 ;
  assign n1323 = n1302 ^ n1298 ;
  assign n1326 = n1322 & n1323 ;
  assign n1320 = n1299 ^ n1295 ;
  assign n1321 = n1300 ^ n1296 ;
  assign n1325 = n1320 & n1321 ;
  assign n1330 = n1326 ^ n1325 ;
  assign n1334 = n1332 ^ n1330 ;
  assign n1335 = n1334 ^ n1319 ;
  assign n1346 = n1340 ^ n1335 ;
  assign n1304 = n1294 ^ n1289 ;
  assign n1347 = n1346 ^ n1304 ;
  assign n1203 = n1182 ^ n1178 ;
  assign n1204 = n1183 ^ n1179 ;
  assign n1207 = n1203 & n1204 ;
  assign n1201 = n1180 ^ n1176 ;
  assign n1202 = n1181 ^ n1177 ;
  assign n1206 = n1201 & n1202 ;
  assign n1211 = n1207 ^ n1206 ;
  assign n1215 = n1213 ^ n1211 ;
  assign n1216 = n1215 ^ n1200 ;
  assign n1227 = n1221 ^ n1216 ;
  assign n1185 = n1175 ^ n1170 ;
  assign n1228 = n1227 ^ n1185 ;
  assign n1498 = n1347 ^ n1228 ;
  assign n1544 = n1522 ^ n1498 ;
  assign n1545 = n1544 ^ n1062 ;
  assign n4295 = n2852 ^ n1545 ;
  assign n12806 = n8407 ^ n4295 ;
  assign n6746 = n6741 ^ n6739 ;
  assign n6747 = n6742 ^ n6740 ;
  assign n6748 = n6746 & n6747 ;
  assign n6750 = n6748 ^ n6744 ;
  assign n6755 = n6752 ^ n6750 ;
  assign n6743 = n6738 ^ n6737 ;
  assign n6756 = n6755 ^ n6743 ;
  assign n6767 = n6760 ^ n6756 ;
  assign n6722 = n6713 ^ n6711 ;
  assign n6724 = n6722 ^ n6709 ;
  assign n6768 = n6767 ^ n6724 ;
  assign n6627 = n6622 ^ n6620 ;
  assign n6628 = n6623 ^ n6621 ;
  assign n6629 = n6627 & n6628 ;
  assign n6631 = n6629 ^ n6625 ;
  assign n6636 = n6633 ^ n6631 ;
  assign n6624 = n6619 ^ n6618 ;
  assign n6637 = n6636 ^ n6624 ;
  assign n6648 = n6641 ^ n6637 ;
  assign n6603 = n6594 ^ n6592 ;
  assign n6605 = n6603 ^ n6590 ;
  assign n6649 = n6648 ^ n6605 ;
  assign n6918 = n6768 ^ n6649 ;
  assign n6965 = n6942 ^ n6918 ;
  assign n6966 = n6965 ^ n6483 ;
  assign n5439 = n5434 ^ n5432 ;
  assign n5440 = n5435 ^ n5433 ;
  assign n5441 = n5439 & n5440 ;
  assign n5443 = n5441 ^ n5437 ;
  assign n5448 = n5445 ^ n5443 ;
  assign n5436 = n5431 ^ n5430 ;
  assign n5449 = n5448 ^ n5436 ;
  assign n5460 = n5453 ^ n5449 ;
  assign n5415 = n5406 ^ n5404 ;
  assign n5417 = n5415 ^ n5402 ;
  assign n5461 = n5460 ^ n5417 ;
  assign n5320 = n5315 ^ n5313 ;
  assign n5321 = n5316 ^ n5314 ;
  assign n5322 = n5320 & n5321 ;
  assign n5324 = n5322 ^ n5318 ;
  assign n5329 = n5326 ^ n5324 ;
  assign n5317 = n5312 ^ n5311 ;
  assign n5330 = n5329 ^ n5317 ;
  assign n5341 = n5334 ^ n5330 ;
  assign n5296 = n5287 ^ n5285 ;
  assign n5298 = n5296 ^ n5283 ;
  assign n5342 = n5341 ^ n5298 ;
  assign n5611 = n5461 ^ n5342 ;
  assign n5658 = n5635 ^ n5611 ;
  assign n5659 = n5658 ^ n5176 ;
  assign n8408 = n6966 ^ n5659 ;
  assign n2634 = n2629 ^ n2627 ;
  assign n2635 = n2630 ^ n2628 ;
  assign n2636 = n2634 & n2635 ;
  assign n2638 = n2636 ^ n2632 ;
  assign n2643 = n2640 ^ n2638 ;
  assign n2631 = n2626 ^ n2625 ;
  assign n2644 = n2643 ^ n2631 ;
  assign n2655 = n2648 ^ n2644 ;
  assign n2610 = n2601 ^ n2599 ;
  assign n2612 = n2610 ^ n2597 ;
  assign n2656 = n2655 ^ n2612 ;
  assign n2515 = n2510 ^ n2508 ;
  assign n2516 = n2511 ^ n2509 ;
  assign n2517 = n2515 & n2516 ;
  assign n2519 = n2517 ^ n2513 ;
  assign n2524 = n2521 ^ n2519 ;
  assign n2512 = n2507 ^ n2506 ;
  assign n2525 = n2524 ^ n2512 ;
  assign n2536 = n2529 ^ n2525 ;
  assign n2491 = n2482 ^ n2480 ;
  assign n2493 = n2491 ^ n2478 ;
  assign n2537 = n2536 ^ n2493 ;
  assign n2806 = n2656 ^ n2537 ;
  assign n2853 = n2830 ^ n2806 ;
  assign n2854 = n2853 ^ n2371 ;
  assign n1327 = n1322 ^ n1320 ;
  assign n1328 = n1323 ^ n1321 ;
  assign n1329 = n1327 & n1328 ;
  assign n1331 = n1329 ^ n1325 ;
  assign n1336 = n1333 ^ n1331 ;
  assign n1324 = n1319 ^ n1318 ;
  assign n1337 = n1336 ^ n1324 ;
  assign n1348 = n1341 ^ n1337 ;
  assign n1303 = n1294 ^ n1292 ;
  assign n1305 = n1303 ^ n1290 ;
  assign n1349 = n1348 ^ n1305 ;
  assign n1208 = n1203 ^ n1201 ;
  assign n1209 = n1204 ^ n1202 ;
  assign n1210 = n1208 & n1209 ;
  assign n1212 = n1210 ^ n1206 ;
  assign n1217 = n1214 ^ n1212 ;
  assign n1205 = n1200 ^ n1199 ;
  assign n1218 = n1217 ^ n1205 ;
  assign n1229 = n1222 ^ n1218 ;
  assign n1184 = n1175 ^ n1173 ;
  assign n1186 = n1184 ^ n1171 ;
  assign n1230 = n1229 ^ n1186 ;
  assign n1499 = n1349 ^ n1230 ;
  assign n1546 = n1523 ^ n1499 ;
  assign n1547 = n1546 ^ n1064 ;
  assign n4296 = n2854 ^ n1547 ;
  assign n12807 = n8408 ^ n4296 ;
  assign n6783 = n6514 ^ n6498 ;
  assign n6784 = n6515 ^ n6499 ;
  assign n6832 = n6783 & n6784 ;
  assign n6781 = n6512 ^ n6496 ;
  assign n6782 = n6513 ^ n6497 ;
  assign n6831 = n6781 & n6782 ;
  assign n6836 = n6832 ^ n6831 ;
  assign n6779 = n6510 ^ n6494 ;
  assign n6780 = n6511 ^ n6495 ;
  assign n6825 = n6779 & n6780 ;
  assign n6777 = n6508 ^ n6492 ;
  assign n6778 = n6509 ^ n6493 ;
  assign n6824 = n6777 & n6778 ;
  assign n6829 = n6825 ^ n6824 ;
  assign n6850 = n6836 ^ n6829 ;
  assign n6775 = n6506 ^ n6490 ;
  assign n6776 = n6507 ^ n6491 ;
  assign n6800 = n6775 & n6776 ;
  assign n6773 = n6504 ^ n6488 ;
  assign n6774 = n6505 ^ n6489 ;
  assign n6799 = n6773 & n6774 ;
  assign n6804 = n6800 ^ n6799 ;
  assign n6771 = n6502 ^ n6486 ;
  assign n6772 = n6503 ^ n6487 ;
  assign n6793 = n6771 & n6772 ;
  assign n6769 = n6500 ^ n6484 ;
  assign n6770 = n6501 ^ n6485 ;
  assign n6792 = n6769 & n6770 ;
  assign n6797 = n6793 ^ n6792 ;
  assign n6818 = n6804 ^ n6797 ;
  assign n6899 = n6850 ^ n6818 ;
  assign n6919 = n6911 ^ n6899 ;
  assign n6920 = n6919 ^ n6762 ;
  assign n6967 = n6943 ^ n6920 ;
  assign n6523 = n6477 ^ n6460 ;
  assign n6968 = n6967 ^ n6523 ;
  assign n5476 = n5207 ^ n5191 ;
  assign n5477 = n5208 ^ n5192 ;
  assign n5525 = n5476 & n5477 ;
  assign n5474 = n5205 ^ n5189 ;
  assign n5475 = n5206 ^ n5190 ;
  assign n5524 = n5474 & n5475 ;
  assign n5529 = n5525 ^ n5524 ;
  assign n5472 = n5203 ^ n5187 ;
  assign n5473 = n5204 ^ n5188 ;
  assign n5518 = n5472 & n5473 ;
  assign n5470 = n5201 ^ n5185 ;
  assign n5471 = n5202 ^ n5186 ;
  assign n5517 = n5470 & n5471 ;
  assign n5522 = n5518 ^ n5517 ;
  assign n5543 = n5529 ^ n5522 ;
  assign n5468 = n5199 ^ n5183 ;
  assign n5469 = n5200 ^ n5184 ;
  assign n5493 = n5468 & n5469 ;
  assign n5466 = n5197 ^ n5181 ;
  assign n5467 = n5198 ^ n5182 ;
  assign n5492 = n5466 & n5467 ;
  assign n5497 = n5493 ^ n5492 ;
  assign n5464 = n5195 ^ n5179 ;
  assign n5465 = n5196 ^ n5180 ;
  assign n5486 = n5464 & n5465 ;
  assign n5462 = n5193 ^ n5177 ;
  assign n5463 = n5194 ^ n5178 ;
  assign n5485 = n5462 & n5463 ;
  assign n5490 = n5486 ^ n5485 ;
  assign n5511 = n5497 ^ n5490 ;
  assign n5592 = n5543 ^ n5511 ;
  assign n5612 = n5604 ^ n5592 ;
  assign n5613 = n5612 ^ n5455 ;
  assign n5660 = n5636 ^ n5613 ;
  assign n5216 = n5170 ^ n5153 ;
  assign n5661 = n5660 ^ n5216 ;
  assign n8409 = n6968 ^ n5661 ;
  assign n2671 = n2402 ^ n2386 ;
  assign n2672 = n2403 ^ n2387 ;
  assign n2720 = n2671 & n2672 ;
  assign n2669 = n2400 ^ n2384 ;
  assign n2670 = n2401 ^ n2385 ;
  assign n2719 = n2669 & n2670 ;
  assign n2724 = n2720 ^ n2719 ;
  assign n2667 = n2398 ^ n2382 ;
  assign n2668 = n2399 ^ n2383 ;
  assign n2713 = n2667 & n2668 ;
  assign n2665 = n2396 ^ n2380 ;
  assign n2666 = n2397 ^ n2381 ;
  assign n2712 = n2665 & n2666 ;
  assign n2717 = n2713 ^ n2712 ;
  assign n2738 = n2724 ^ n2717 ;
  assign n2663 = n2394 ^ n2378 ;
  assign n2664 = n2395 ^ n2379 ;
  assign n2688 = n2663 & n2664 ;
  assign n2661 = n2392 ^ n2376 ;
  assign n2662 = n2393 ^ n2377 ;
  assign n2687 = n2661 & n2662 ;
  assign n2692 = n2688 ^ n2687 ;
  assign n2659 = n2390 ^ n2374 ;
  assign n2660 = n2391 ^ n2375 ;
  assign n2681 = n2659 & n2660 ;
  assign n2657 = n2388 ^ n2372 ;
  assign n2658 = n2389 ^ n2373 ;
  assign n2680 = n2657 & n2658 ;
  assign n2685 = n2681 ^ n2680 ;
  assign n2706 = n2692 ^ n2685 ;
  assign n2787 = n2738 ^ n2706 ;
  assign n2807 = n2799 ^ n2787 ;
  assign n2808 = n2807 ^ n2650 ;
  assign n2855 = n2831 ^ n2808 ;
  assign n2411 = n2365 ^ n2348 ;
  assign n2856 = n2855 ^ n2411 ;
  assign n1364 = n1095 ^ n1079 ;
  assign n1365 = n1096 ^ n1080 ;
  assign n1413 = n1364 & n1365 ;
  assign n1362 = n1093 ^ n1077 ;
  assign n1363 = n1094 ^ n1078 ;
  assign n1412 = n1362 & n1363 ;
  assign n1417 = n1413 ^ n1412 ;
  assign n1360 = n1091 ^ n1075 ;
  assign n1361 = n1092 ^ n1076 ;
  assign n1406 = n1360 & n1361 ;
  assign n1358 = n1089 ^ n1073 ;
  assign n1359 = n1090 ^ n1074 ;
  assign n1405 = n1358 & n1359 ;
  assign n1410 = n1406 ^ n1405 ;
  assign n1431 = n1417 ^ n1410 ;
  assign n1356 = n1087 ^ n1071 ;
  assign n1357 = n1088 ^ n1072 ;
  assign n1381 = n1356 & n1357 ;
  assign n1354 = n1085 ^ n1069 ;
  assign n1355 = n1086 ^ n1070 ;
  assign n1380 = n1354 & n1355 ;
  assign n1385 = n1381 ^ n1380 ;
  assign n1352 = n1083 ^ n1067 ;
  assign n1353 = n1084 ^ n1068 ;
  assign n1374 = n1352 & n1353 ;
  assign n1350 = n1081 ^ n1065 ;
  assign n1351 = n1082 ^ n1066 ;
  assign n1373 = n1350 & n1351 ;
  assign n1378 = n1374 ^ n1373 ;
  assign n1399 = n1385 ^ n1378 ;
  assign n1480 = n1431 ^ n1399 ;
  assign n1500 = n1492 ^ n1480 ;
  assign n1501 = n1500 ^ n1343 ;
  assign n1548 = n1524 ^ n1501 ;
  assign n1104 = n1058 ^ n1041 ;
  assign n1549 = n1548 ^ n1104 ;
  assign n4297 = n2856 ^ n1549 ;
  assign n12808 = n8409 ^ n4297 ;
  assign n6833 = n6783 ^ n6781 ;
  assign n6834 = n6784 ^ n6782 ;
  assign n6835 = n6833 & n6834 ;
  assign n6837 = n6835 ^ n6831 ;
  assign n6826 = n6779 ^ n6777 ;
  assign n6827 = n6780 ^ n6778 ;
  assign n6828 = n6826 & n6827 ;
  assign n6830 = n6828 ^ n6824 ;
  assign n6851 = n6837 ^ n6830 ;
  assign n6801 = n6775 ^ n6773 ;
  assign n6802 = n6776 ^ n6774 ;
  assign n6803 = n6801 & n6802 ;
  assign n6805 = n6803 ^ n6799 ;
  assign n6794 = n6771 ^ n6769 ;
  assign n6795 = n6772 ^ n6770 ;
  assign n6796 = n6794 & n6795 ;
  assign n6798 = n6796 ^ n6792 ;
  assign n6819 = n6805 ^ n6798 ;
  assign n6900 = n6851 ^ n6819 ;
  assign n6921 = n6912 ^ n6900 ;
  assign n6922 = n6921 ^ n6764 ;
  assign n6969 = n6944 ^ n6922 ;
  assign n6524 = n6479 ^ n6461 ;
  assign n6970 = n6969 ^ n6524 ;
  assign n5526 = n5476 ^ n5474 ;
  assign n5527 = n5477 ^ n5475 ;
  assign n5528 = n5526 & n5527 ;
  assign n5530 = n5528 ^ n5524 ;
  assign n5519 = n5472 ^ n5470 ;
  assign n5520 = n5473 ^ n5471 ;
  assign n5521 = n5519 & n5520 ;
  assign n5523 = n5521 ^ n5517 ;
  assign n5544 = n5530 ^ n5523 ;
  assign n5494 = n5468 ^ n5466 ;
  assign n5495 = n5469 ^ n5467 ;
  assign n5496 = n5494 & n5495 ;
  assign n5498 = n5496 ^ n5492 ;
  assign n5487 = n5464 ^ n5462 ;
  assign n5488 = n5465 ^ n5463 ;
  assign n5489 = n5487 & n5488 ;
  assign n5491 = n5489 ^ n5485 ;
  assign n5512 = n5498 ^ n5491 ;
  assign n5593 = n5544 ^ n5512 ;
  assign n5614 = n5605 ^ n5593 ;
  assign n5615 = n5614 ^ n5457 ;
  assign n5662 = n5637 ^ n5615 ;
  assign n5217 = n5172 ^ n5154 ;
  assign n5663 = n5662 ^ n5217 ;
  assign n8410 = n6970 ^ n5663 ;
  assign n2721 = n2671 ^ n2669 ;
  assign n2722 = n2672 ^ n2670 ;
  assign n2723 = n2721 & n2722 ;
  assign n2725 = n2723 ^ n2719 ;
  assign n2714 = n2667 ^ n2665 ;
  assign n2715 = n2668 ^ n2666 ;
  assign n2716 = n2714 & n2715 ;
  assign n2718 = n2716 ^ n2712 ;
  assign n2739 = n2725 ^ n2718 ;
  assign n2689 = n2663 ^ n2661 ;
  assign n2690 = n2664 ^ n2662 ;
  assign n2691 = n2689 & n2690 ;
  assign n2693 = n2691 ^ n2687 ;
  assign n2682 = n2659 ^ n2657 ;
  assign n2683 = n2660 ^ n2658 ;
  assign n2684 = n2682 & n2683 ;
  assign n2686 = n2684 ^ n2680 ;
  assign n2707 = n2693 ^ n2686 ;
  assign n2788 = n2739 ^ n2707 ;
  assign n2809 = n2800 ^ n2788 ;
  assign n2810 = n2809 ^ n2652 ;
  assign n2857 = n2832 ^ n2810 ;
  assign n2412 = n2367 ^ n2349 ;
  assign n2858 = n2857 ^ n2412 ;
  assign n1414 = n1364 ^ n1362 ;
  assign n1415 = n1365 ^ n1363 ;
  assign n1416 = n1414 & n1415 ;
  assign n1418 = n1416 ^ n1412 ;
  assign n1407 = n1360 ^ n1358 ;
  assign n1408 = n1361 ^ n1359 ;
  assign n1409 = n1407 & n1408 ;
  assign n1411 = n1409 ^ n1405 ;
  assign n1432 = n1418 ^ n1411 ;
  assign n1382 = n1356 ^ n1354 ;
  assign n1383 = n1357 ^ n1355 ;
  assign n1384 = n1382 & n1383 ;
  assign n1386 = n1384 ^ n1380 ;
  assign n1375 = n1352 ^ n1350 ;
  assign n1376 = n1353 ^ n1351 ;
  assign n1377 = n1375 & n1376 ;
  assign n1379 = n1377 ^ n1373 ;
  assign n1400 = n1386 ^ n1379 ;
  assign n1481 = n1432 ^ n1400 ;
  assign n1502 = n1493 ^ n1481 ;
  assign n1503 = n1502 ^ n1345 ;
  assign n1550 = n1525 ^ n1503 ;
  assign n1105 = n1060 ^ n1042 ;
  assign n1551 = n1550 ^ n1105 ;
  assign n4298 = n2858 ^ n1551 ;
  assign n12809 = n8410 ^ n4298 ;
  assign n6840 = n6783 ^ n6779 ;
  assign n6841 = n6784 ^ n6780 ;
  assign n6844 = n6840 & n6841 ;
  assign n6838 = n6781 ^ n6777 ;
  assign n6839 = n6782 ^ n6778 ;
  assign n6843 = n6838 & n6839 ;
  assign n6848 = n6844 ^ n6843 ;
  assign n6852 = n6850 ^ n6848 ;
  assign n6853 = n6852 ^ n6837 ;
  assign n6808 = n6775 ^ n6771 ;
  assign n6809 = n6776 ^ n6772 ;
  assign n6812 = n6808 & n6809 ;
  assign n6806 = n6773 ^ n6769 ;
  assign n6807 = n6774 ^ n6770 ;
  assign n6811 = n6806 & n6807 ;
  assign n6816 = n6812 ^ n6811 ;
  assign n6820 = n6818 ^ n6816 ;
  assign n6821 = n6820 ^ n6805 ;
  assign n6901 = n6853 ^ n6821 ;
  assign n6923 = n6913 ^ n6901 ;
  assign n6924 = n6923 ^ n6766 ;
  assign n6971 = n6945 ^ n6924 ;
  assign n6525 = n6481 ^ n6462 ;
  assign n6972 = n6971 ^ n6525 ;
  assign n5533 = n5476 ^ n5472 ;
  assign n5534 = n5477 ^ n5473 ;
  assign n5537 = n5533 & n5534 ;
  assign n5531 = n5474 ^ n5470 ;
  assign n5532 = n5475 ^ n5471 ;
  assign n5536 = n5531 & n5532 ;
  assign n5541 = n5537 ^ n5536 ;
  assign n5545 = n5543 ^ n5541 ;
  assign n5546 = n5545 ^ n5530 ;
  assign n5501 = n5468 ^ n5464 ;
  assign n5502 = n5469 ^ n5465 ;
  assign n5505 = n5501 & n5502 ;
  assign n5499 = n5466 ^ n5462 ;
  assign n5500 = n5467 ^ n5463 ;
  assign n5504 = n5499 & n5500 ;
  assign n5509 = n5505 ^ n5504 ;
  assign n5513 = n5511 ^ n5509 ;
  assign n5514 = n5513 ^ n5498 ;
  assign n5594 = n5546 ^ n5514 ;
  assign n5616 = n5606 ^ n5594 ;
  assign n5617 = n5616 ^ n5459 ;
  assign n5664 = n5638 ^ n5617 ;
  assign n5218 = n5174 ^ n5155 ;
  assign n5665 = n5664 ^ n5218 ;
  assign n8411 = n6972 ^ n5665 ;
  assign n2728 = n2671 ^ n2667 ;
  assign n2729 = n2672 ^ n2668 ;
  assign n2732 = n2728 & n2729 ;
  assign n2726 = n2669 ^ n2665 ;
  assign n2727 = n2670 ^ n2666 ;
  assign n2731 = n2726 & n2727 ;
  assign n2736 = n2732 ^ n2731 ;
  assign n2740 = n2738 ^ n2736 ;
  assign n2741 = n2740 ^ n2725 ;
  assign n2696 = n2663 ^ n2659 ;
  assign n2697 = n2664 ^ n2660 ;
  assign n2700 = n2696 & n2697 ;
  assign n2694 = n2661 ^ n2657 ;
  assign n2695 = n2662 ^ n2658 ;
  assign n2699 = n2694 & n2695 ;
  assign n2704 = n2700 ^ n2699 ;
  assign n2708 = n2706 ^ n2704 ;
  assign n2709 = n2708 ^ n2693 ;
  assign n2789 = n2741 ^ n2709 ;
  assign n2811 = n2801 ^ n2789 ;
  assign n2812 = n2811 ^ n2654 ;
  assign n2859 = n2833 ^ n2812 ;
  assign n2413 = n2369 ^ n2350 ;
  assign n2860 = n2859 ^ n2413 ;
  assign n1421 = n1364 ^ n1360 ;
  assign n1422 = n1365 ^ n1361 ;
  assign n1425 = n1421 & n1422 ;
  assign n1419 = n1362 ^ n1358 ;
  assign n1420 = n1363 ^ n1359 ;
  assign n1424 = n1419 & n1420 ;
  assign n1429 = n1425 ^ n1424 ;
  assign n1433 = n1431 ^ n1429 ;
  assign n1434 = n1433 ^ n1418 ;
  assign n1389 = n1356 ^ n1352 ;
  assign n1390 = n1357 ^ n1353 ;
  assign n1393 = n1389 & n1390 ;
  assign n1387 = n1354 ^ n1350 ;
  assign n1388 = n1355 ^ n1351 ;
  assign n1392 = n1387 & n1388 ;
  assign n1397 = n1393 ^ n1392 ;
  assign n1401 = n1399 ^ n1397 ;
  assign n1402 = n1401 ^ n1386 ;
  assign n1482 = n1434 ^ n1402 ;
  assign n1504 = n1494 ^ n1482 ;
  assign n1505 = n1504 ^ n1347 ;
  assign n1552 = n1526 ^ n1505 ;
  assign n1106 = n1062 ^ n1043 ;
  assign n1553 = n1552 ^ n1106 ;
  assign n4299 = n2860 ^ n1553 ;
  assign n12810 = n8411 ^ n4299 ;
  assign n6845 = n6840 ^ n6838 ;
  assign n6846 = n6841 ^ n6839 ;
  assign n6847 = n6845 & n6846 ;
  assign n6849 = n6847 ^ n6843 ;
  assign n6854 = n6851 ^ n6849 ;
  assign n6842 = n6837 ^ n6836 ;
  assign n6855 = n6854 ^ n6842 ;
  assign n6813 = n6808 ^ n6806 ;
  assign n6814 = n6809 ^ n6807 ;
  assign n6815 = n6813 & n6814 ;
  assign n6817 = n6815 ^ n6811 ;
  assign n6822 = n6819 ^ n6817 ;
  assign n6810 = n6805 ^ n6804 ;
  assign n6823 = n6822 ^ n6810 ;
  assign n6902 = n6855 ^ n6823 ;
  assign n6925 = n6914 ^ n6902 ;
  assign n6926 = n6925 ^ n6768 ;
  assign n6973 = n6946 ^ n6926 ;
  assign n6526 = n6483 ^ n6463 ;
  assign n6974 = n6973 ^ n6526 ;
  assign n5538 = n5533 ^ n5531 ;
  assign n5539 = n5534 ^ n5532 ;
  assign n5540 = n5538 & n5539 ;
  assign n5542 = n5540 ^ n5536 ;
  assign n5547 = n5544 ^ n5542 ;
  assign n5535 = n5530 ^ n5529 ;
  assign n5548 = n5547 ^ n5535 ;
  assign n5506 = n5501 ^ n5499 ;
  assign n5507 = n5502 ^ n5500 ;
  assign n5508 = n5506 & n5507 ;
  assign n5510 = n5508 ^ n5504 ;
  assign n5515 = n5512 ^ n5510 ;
  assign n5503 = n5498 ^ n5497 ;
  assign n5516 = n5515 ^ n5503 ;
  assign n5595 = n5548 ^ n5516 ;
  assign n5618 = n5607 ^ n5595 ;
  assign n5619 = n5618 ^ n5461 ;
  assign n5666 = n5639 ^ n5619 ;
  assign n5219 = n5176 ^ n5156 ;
  assign n5667 = n5666 ^ n5219 ;
  assign n8412 = n6974 ^ n5667 ;
  assign n2733 = n2728 ^ n2726 ;
  assign n2734 = n2729 ^ n2727 ;
  assign n2735 = n2733 & n2734 ;
  assign n2737 = n2735 ^ n2731 ;
  assign n2742 = n2739 ^ n2737 ;
  assign n2730 = n2725 ^ n2724 ;
  assign n2743 = n2742 ^ n2730 ;
  assign n2701 = n2696 ^ n2694 ;
  assign n2702 = n2697 ^ n2695 ;
  assign n2703 = n2701 & n2702 ;
  assign n2705 = n2703 ^ n2699 ;
  assign n2710 = n2707 ^ n2705 ;
  assign n2698 = n2693 ^ n2692 ;
  assign n2711 = n2710 ^ n2698 ;
  assign n2790 = n2743 ^ n2711 ;
  assign n2813 = n2802 ^ n2790 ;
  assign n2814 = n2813 ^ n2656 ;
  assign n2861 = n2834 ^ n2814 ;
  assign n2414 = n2371 ^ n2351 ;
  assign n2862 = n2861 ^ n2414 ;
  assign n1426 = n1421 ^ n1419 ;
  assign n1427 = n1422 ^ n1420 ;
  assign n1428 = n1426 & n1427 ;
  assign n1430 = n1428 ^ n1424 ;
  assign n1435 = n1432 ^ n1430 ;
  assign n1423 = n1418 ^ n1417 ;
  assign n1436 = n1435 ^ n1423 ;
  assign n1394 = n1389 ^ n1387 ;
  assign n1395 = n1390 ^ n1388 ;
  assign n1396 = n1394 & n1395 ;
  assign n1398 = n1396 ^ n1392 ;
  assign n1403 = n1400 ^ n1398 ;
  assign n1391 = n1386 ^ n1385 ;
  assign n1404 = n1403 ^ n1391 ;
  assign n1483 = n1436 ^ n1404 ;
  assign n1506 = n1495 ^ n1483 ;
  assign n1507 = n1506 ^ n1349 ;
  assign n1554 = n1527 ^ n1507 ;
  assign n1107 = n1064 ^ n1044 ;
  assign n1555 = n1554 ^ n1107 ;
  assign n4300 = n2862 ^ n1555 ;
  assign n12811 = n8412 ^ n4300 ;
  assign n6862 = n6783 ^ n6775 ;
  assign n6863 = n6784 ^ n6776 ;
  assign n6875 = n6862 & n6863 ;
  assign n6860 = n6781 ^ n6773 ;
  assign n6861 = n6782 ^ n6774 ;
  assign n6874 = n6860 & n6861 ;
  assign n6879 = n6875 ^ n6874 ;
  assign n6858 = n6779 ^ n6771 ;
  assign n6859 = n6780 ^ n6772 ;
  assign n6868 = n6858 & n6859 ;
  assign n6856 = n6777 ^ n6769 ;
  assign n6857 = n6778 ^ n6770 ;
  assign n6867 = n6856 & n6857 ;
  assign n6872 = n6868 ^ n6867 ;
  assign n6893 = n6879 ^ n6872 ;
  assign n6903 = n6899 ^ n6893 ;
  assign n6904 = n6903 ^ n6853 ;
  assign n6927 = n6915 ^ n6904 ;
  assign n6788 = n6766 ^ n6757 ;
  assign n6928 = n6927 ^ n6788 ;
  assign n6975 = n6947 ^ n6928 ;
  assign n6519 = n6481 ^ n6469 ;
  assign n6527 = n6519 ^ n6464 ;
  assign n6976 = n6975 ^ n6527 ;
  assign n5555 = n5476 ^ n5468 ;
  assign n5556 = n5477 ^ n5469 ;
  assign n5568 = n5555 & n5556 ;
  assign n5553 = n5474 ^ n5466 ;
  assign n5554 = n5475 ^ n5467 ;
  assign n5567 = n5553 & n5554 ;
  assign n5572 = n5568 ^ n5567 ;
  assign n5551 = n5472 ^ n5464 ;
  assign n5552 = n5473 ^ n5465 ;
  assign n5561 = n5551 & n5552 ;
  assign n5549 = n5470 ^ n5462 ;
  assign n5550 = n5471 ^ n5463 ;
  assign n5560 = n5549 & n5550 ;
  assign n5565 = n5561 ^ n5560 ;
  assign n5586 = n5572 ^ n5565 ;
  assign n5596 = n5592 ^ n5586 ;
  assign n5597 = n5596 ^ n5546 ;
  assign n5620 = n5608 ^ n5597 ;
  assign n5481 = n5459 ^ n5450 ;
  assign n5621 = n5620 ^ n5481 ;
  assign n5668 = n5640 ^ n5621 ;
  assign n5212 = n5174 ^ n5162 ;
  assign n5220 = n5212 ^ n5157 ;
  assign n5669 = n5668 ^ n5220 ;
  assign n8413 = n6976 ^ n5669 ;
  assign n2750 = n2671 ^ n2663 ;
  assign n2751 = n2672 ^ n2664 ;
  assign n2763 = n2750 & n2751 ;
  assign n2748 = n2669 ^ n2661 ;
  assign n2749 = n2670 ^ n2662 ;
  assign n2762 = n2748 & n2749 ;
  assign n2767 = n2763 ^ n2762 ;
  assign n2746 = n2667 ^ n2659 ;
  assign n2747 = n2668 ^ n2660 ;
  assign n2756 = n2746 & n2747 ;
  assign n2744 = n2665 ^ n2657 ;
  assign n2745 = n2666 ^ n2658 ;
  assign n2755 = n2744 & n2745 ;
  assign n2760 = n2756 ^ n2755 ;
  assign n2781 = n2767 ^ n2760 ;
  assign n2791 = n2787 ^ n2781 ;
  assign n2792 = n2791 ^ n2741 ;
  assign n2815 = n2803 ^ n2792 ;
  assign n2676 = n2654 ^ n2645 ;
  assign n2816 = n2815 ^ n2676 ;
  assign n2863 = n2835 ^ n2816 ;
  assign n2407 = n2369 ^ n2357 ;
  assign n2415 = n2407 ^ n2352 ;
  assign n2864 = n2863 ^ n2415 ;
  assign n1443 = n1364 ^ n1356 ;
  assign n1444 = n1365 ^ n1357 ;
  assign n1456 = n1443 & n1444 ;
  assign n1441 = n1362 ^ n1354 ;
  assign n1442 = n1363 ^ n1355 ;
  assign n1455 = n1441 & n1442 ;
  assign n1460 = n1456 ^ n1455 ;
  assign n1439 = n1360 ^ n1352 ;
  assign n1440 = n1361 ^ n1353 ;
  assign n1449 = n1439 & n1440 ;
  assign n1437 = n1358 ^ n1350 ;
  assign n1438 = n1359 ^ n1351 ;
  assign n1448 = n1437 & n1438 ;
  assign n1453 = n1449 ^ n1448 ;
  assign n1474 = n1460 ^ n1453 ;
  assign n1484 = n1480 ^ n1474 ;
  assign n1485 = n1484 ^ n1434 ;
  assign n1508 = n1496 ^ n1485 ;
  assign n1369 = n1347 ^ n1338 ;
  assign n1509 = n1508 ^ n1369 ;
  assign n1556 = n1528 ^ n1509 ;
  assign n1100 = n1062 ^ n1050 ;
  assign n1108 = n1100 ^ n1045 ;
  assign n1557 = n1556 ^ n1108 ;
  assign n4301 = n2864 ^ n1557 ;
  assign n12812 = n8413 ^ n4301 ;
  assign n6876 = n6862 ^ n6860 ;
  assign n6877 = n6863 ^ n6861 ;
  assign n6878 = n6876 & n6877 ;
  assign n6880 = n6878 ^ n6874 ;
  assign n6869 = n6858 ^ n6856 ;
  assign n6870 = n6859 ^ n6857 ;
  assign n6871 = n6869 & n6870 ;
  assign n6873 = n6871 ^ n6867 ;
  assign n6894 = n6880 ^ n6873 ;
  assign n6905 = n6900 ^ n6894 ;
  assign n6906 = n6905 ^ n6855 ;
  assign n6929 = n6916 ^ n6906 ;
  assign n6789 = n6768 ^ n6758 ;
  assign n6930 = n6929 ^ n6789 ;
  assign n6977 = n6948 ^ n6930 ;
  assign n6520 = n6483 ^ n6471 ;
  assign n6528 = n6520 ^ n6465 ;
  assign n6978 = n6977 ^ n6528 ;
  assign n5569 = n5555 ^ n5553 ;
  assign n5570 = n5556 ^ n5554 ;
  assign n5571 = n5569 & n5570 ;
  assign n5573 = n5571 ^ n5567 ;
  assign n5562 = n5551 ^ n5549 ;
  assign n5563 = n5552 ^ n5550 ;
  assign n5564 = n5562 & n5563 ;
  assign n5566 = n5564 ^ n5560 ;
  assign n5587 = n5573 ^ n5566 ;
  assign n5598 = n5593 ^ n5587 ;
  assign n5599 = n5598 ^ n5548 ;
  assign n5622 = n5609 ^ n5599 ;
  assign n5482 = n5461 ^ n5451 ;
  assign n5623 = n5622 ^ n5482 ;
  assign n5670 = n5641 ^ n5623 ;
  assign n5213 = n5176 ^ n5164 ;
  assign n5221 = n5213 ^ n5158 ;
  assign n5671 = n5670 ^ n5221 ;
  assign n8414 = n6978 ^ n5671 ;
  assign n2764 = n2750 ^ n2748 ;
  assign n2765 = n2751 ^ n2749 ;
  assign n2766 = n2764 & n2765 ;
  assign n2768 = n2766 ^ n2762 ;
  assign n2757 = n2746 ^ n2744 ;
  assign n2758 = n2747 ^ n2745 ;
  assign n2759 = n2757 & n2758 ;
  assign n2761 = n2759 ^ n2755 ;
  assign n2782 = n2768 ^ n2761 ;
  assign n2793 = n2788 ^ n2782 ;
  assign n2794 = n2793 ^ n2743 ;
  assign n2817 = n2804 ^ n2794 ;
  assign n2677 = n2656 ^ n2646 ;
  assign n2818 = n2817 ^ n2677 ;
  assign n2865 = n2836 ^ n2818 ;
  assign n2408 = n2371 ^ n2359 ;
  assign n2416 = n2408 ^ n2353 ;
  assign n2866 = n2865 ^ n2416 ;
  assign n1457 = n1443 ^ n1441 ;
  assign n1458 = n1444 ^ n1442 ;
  assign n1459 = n1457 & n1458 ;
  assign n1461 = n1459 ^ n1455 ;
  assign n1450 = n1439 ^ n1437 ;
  assign n1451 = n1440 ^ n1438 ;
  assign n1452 = n1450 & n1451 ;
  assign n1454 = n1452 ^ n1448 ;
  assign n1475 = n1461 ^ n1454 ;
  assign n1486 = n1481 ^ n1475 ;
  assign n1487 = n1486 ^ n1436 ;
  assign n1510 = n1497 ^ n1487 ;
  assign n1370 = n1349 ^ n1339 ;
  assign n1511 = n1510 ^ n1370 ;
  assign n1558 = n1529 ^ n1511 ;
  assign n1101 = n1064 ^ n1052 ;
  assign n1109 = n1101 ^ n1046 ;
  assign n1559 = n1558 ^ n1109 ;
  assign n4302 = n2866 ^ n1559 ;
  assign n12813 = n8414 ^ n4302 ;
  assign n6883 = n6862 ^ n6858 ;
  assign n6884 = n6863 ^ n6859 ;
  assign n6887 = n6883 & n6884 ;
  assign n6881 = n6860 ^ n6856 ;
  assign n6882 = n6861 ^ n6857 ;
  assign n6886 = n6881 & n6882 ;
  assign n6891 = n6887 ^ n6886 ;
  assign n6895 = n6893 ^ n6891 ;
  assign n6896 = n6895 ^ n6880 ;
  assign n6907 = n6901 ^ n6896 ;
  assign n6865 = n6855 ^ n6850 ;
  assign n6908 = n6907 ^ n6865 ;
  assign n6931 = n6917 ^ n6908 ;
  assign n6786 = n6768 ^ n6762 ;
  assign n6790 = n6786 ^ n6759 ;
  assign n6932 = n6931 ^ n6790 ;
  assign n6979 = n6949 ^ n6932 ;
  assign n6517 = n6483 ^ n6477 ;
  assign n6521 = n6517 ^ n6473 ;
  assign n6529 = n6521 ^ n6466 ;
  assign n6980 = n6979 ^ n6529 ;
  assign n5576 = n5555 ^ n5551 ;
  assign n5577 = n5556 ^ n5552 ;
  assign n5580 = n5576 & n5577 ;
  assign n5574 = n5553 ^ n5549 ;
  assign n5575 = n5554 ^ n5550 ;
  assign n5579 = n5574 & n5575 ;
  assign n5584 = n5580 ^ n5579 ;
  assign n5588 = n5586 ^ n5584 ;
  assign n5589 = n5588 ^ n5573 ;
  assign n5600 = n5594 ^ n5589 ;
  assign n5558 = n5548 ^ n5543 ;
  assign n5601 = n5600 ^ n5558 ;
  assign n5624 = n5610 ^ n5601 ;
  assign n5479 = n5461 ^ n5455 ;
  assign n5483 = n5479 ^ n5452 ;
  assign n5625 = n5624 ^ n5483 ;
  assign n5672 = n5642 ^ n5625 ;
  assign n5210 = n5176 ^ n5170 ;
  assign n5214 = n5210 ^ n5166 ;
  assign n5222 = n5214 ^ n5159 ;
  assign n5673 = n5672 ^ n5222 ;
  assign n8415 = n6980 ^ n5673 ;
  assign n2771 = n2750 ^ n2746 ;
  assign n2772 = n2751 ^ n2747 ;
  assign n2775 = n2771 & n2772 ;
  assign n2769 = n2748 ^ n2744 ;
  assign n2770 = n2749 ^ n2745 ;
  assign n2774 = n2769 & n2770 ;
  assign n2779 = n2775 ^ n2774 ;
  assign n2783 = n2781 ^ n2779 ;
  assign n2784 = n2783 ^ n2768 ;
  assign n2795 = n2789 ^ n2784 ;
  assign n2753 = n2743 ^ n2738 ;
  assign n2796 = n2795 ^ n2753 ;
  assign n2819 = n2805 ^ n2796 ;
  assign n2674 = n2656 ^ n2650 ;
  assign n2678 = n2674 ^ n2647 ;
  assign n2820 = n2819 ^ n2678 ;
  assign n2867 = n2837 ^ n2820 ;
  assign n2405 = n2371 ^ n2365 ;
  assign n2409 = n2405 ^ n2361 ;
  assign n2417 = n2409 ^ n2354 ;
  assign n2868 = n2867 ^ n2417 ;
  assign n1464 = n1443 ^ n1439 ;
  assign n1465 = n1444 ^ n1440 ;
  assign n1468 = n1464 & n1465 ;
  assign n1462 = n1441 ^ n1437 ;
  assign n1463 = n1442 ^ n1438 ;
  assign n1467 = n1462 & n1463 ;
  assign n1472 = n1468 ^ n1467 ;
  assign n1476 = n1474 ^ n1472 ;
  assign n1477 = n1476 ^ n1461 ;
  assign n1488 = n1482 ^ n1477 ;
  assign n1446 = n1436 ^ n1431 ;
  assign n1489 = n1488 ^ n1446 ;
  assign n1512 = n1498 ^ n1489 ;
  assign n1367 = n1349 ^ n1343 ;
  assign n1371 = n1367 ^ n1340 ;
  assign n1513 = n1512 ^ n1371 ;
  assign n1560 = n1530 ^ n1513 ;
  assign n1098 = n1064 ^ n1058 ;
  assign n1102 = n1098 ^ n1054 ;
  assign n1110 = n1102 ^ n1047 ;
  assign n1561 = n1560 ^ n1110 ;
  assign n4303 = n2868 ^ n1561 ;
  assign n12814 = n8415 ^ n4303 ;
  assign n6888 = n6883 ^ n6881 ;
  assign n6889 = n6884 ^ n6882 ;
  assign n6890 = n6888 & n6889 ;
  assign n6892 = n6890 ^ n6886 ;
  assign n6897 = n6894 ^ n6892 ;
  assign n6885 = n6880 ^ n6879 ;
  assign n6898 = n6897 ^ n6885 ;
  assign n6909 = n6902 ^ n6898 ;
  assign n6864 = n6855 ^ n6853 ;
  assign n6866 = n6864 ^ n6851 ;
  assign n6910 = n6909 ^ n6866 ;
  assign n6933 = n6918 ^ n6910 ;
  assign n6785 = n6768 ^ n6766 ;
  assign n6787 = n6785 ^ n6764 ;
  assign n6791 = n6787 ^ n6760 ;
  assign n6934 = n6933 ^ n6791 ;
  assign n6981 = n6950 ^ n6934 ;
  assign n6516 = n6483 ^ n6481 ;
  assign n6518 = n6516 ^ n6479 ;
  assign n6522 = n6518 ^ n6475 ;
  assign n6530 = n6522 ^ n6467 ;
  assign n6982 = n6981 ^ n6530 ;
  assign n5581 = n5576 ^ n5574 ;
  assign n5582 = n5577 ^ n5575 ;
  assign n5583 = n5581 & n5582 ;
  assign n5585 = n5583 ^ n5579 ;
  assign n5590 = n5587 ^ n5585 ;
  assign n5578 = n5573 ^ n5572 ;
  assign n5591 = n5590 ^ n5578 ;
  assign n5602 = n5595 ^ n5591 ;
  assign n5557 = n5548 ^ n5546 ;
  assign n5559 = n5557 ^ n5544 ;
  assign n5603 = n5602 ^ n5559 ;
  assign n5626 = n5611 ^ n5603 ;
  assign n5478 = n5461 ^ n5459 ;
  assign n5480 = n5478 ^ n5457 ;
  assign n5484 = n5480 ^ n5453 ;
  assign n5627 = n5626 ^ n5484 ;
  assign n5674 = n5643 ^ n5627 ;
  assign n5209 = n5176 ^ n5174 ;
  assign n5211 = n5209 ^ n5172 ;
  assign n5215 = n5211 ^ n5168 ;
  assign n5223 = n5215 ^ n5160 ;
  assign n5675 = n5674 ^ n5223 ;
  assign n8416 = n6982 ^ n5675 ;
  assign n2776 = n2771 ^ n2769 ;
  assign n2777 = n2772 ^ n2770 ;
  assign n2778 = n2776 & n2777 ;
  assign n2780 = n2778 ^ n2774 ;
  assign n2785 = n2782 ^ n2780 ;
  assign n2773 = n2768 ^ n2767 ;
  assign n2786 = n2785 ^ n2773 ;
  assign n2797 = n2790 ^ n2786 ;
  assign n2752 = n2743 ^ n2741 ;
  assign n2754 = n2752 ^ n2739 ;
  assign n2798 = n2797 ^ n2754 ;
  assign n2821 = n2806 ^ n2798 ;
  assign n2673 = n2656 ^ n2654 ;
  assign n2675 = n2673 ^ n2652 ;
  assign n2679 = n2675 ^ n2648 ;
  assign n2822 = n2821 ^ n2679 ;
  assign n2869 = n2838 ^ n2822 ;
  assign n2404 = n2371 ^ n2369 ;
  assign n2406 = n2404 ^ n2367 ;
  assign n2410 = n2406 ^ n2363 ;
  assign n2418 = n2410 ^ n2355 ;
  assign n2870 = n2869 ^ n2418 ;
  assign n1469 = n1464 ^ n1462 ;
  assign n1470 = n1465 ^ n1463 ;
  assign n1471 = n1469 & n1470 ;
  assign n1473 = n1471 ^ n1467 ;
  assign n1478 = n1475 ^ n1473 ;
  assign n1466 = n1461 ^ n1460 ;
  assign n1479 = n1478 ^ n1466 ;
  assign n1490 = n1483 ^ n1479 ;
  assign n1445 = n1436 ^ n1434 ;
  assign n1447 = n1445 ^ n1432 ;
  assign n1491 = n1490 ^ n1447 ;
  assign n1514 = n1499 ^ n1491 ;
  assign n1366 = n1349 ^ n1347 ;
  assign n1368 = n1366 ^ n1345 ;
  assign n1372 = n1368 ^ n1341 ;
  assign n1515 = n1514 ^ n1372 ;
  assign n1562 = n1531 ^ n1515 ;
  assign n1097 = n1064 ^ n1062 ;
  assign n1099 = n1097 ^ n1060 ;
  assign n1103 = n1099 ^ n1056 ;
  assign n1111 = n1103 ^ n1048 ;
  assign n1563 = n1562 ^ n1111 ;
  assign n4304 = n2870 ^ n1563 ;
  assign n12815 = n8416 ^ n4304 ;
  assign n7045 = x127 ^ x95 ;
  assign n7046 = x255 ^ x223 ;
  assign n7641 = n7045 & n7046 ;
  assign n7043 = x126 ^ x94 ;
  assign n7044 = x254 ^ x222 ;
  assign n7640 = n7043 & n7044 ;
  assign n7645 = n7641 ^ n7640 ;
  assign n7041 = x125 ^ x93 ;
  assign n7042 = x253 ^ x221 ;
  assign n7634 = n7041 & n7042 ;
  assign n7039 = x124 ^ x92 ;
  assign n7040 = x252 ^ x220 ;
  assign n7633 = n7039 & n7040 ;
  assign n7638 = n7634 ^ n7633 ;
  assign n7659 = n7645 ^ n7638 ;
  assign n7037 = x123 ^ x91 ;
  assign n7038 = x251 ^ x219 ;
  assign n7609 = n7037 & n7038 ;
  assign n7035 = x122 ^ x90 ;
  assign n7036 = x250 ^ x218 ;
  assign n7608 = n7035 & n7036 ;
  assign n7613 = n7609 ^ n7608 ;
  assign n7033 = x121 ^ x89 ;
  assign n7034 = x249 ^ x217 ;
  assign n7602 = n7033 & n7034 ;
  assign n7031 = x120 ^ x88 ;
  assign n7032 = x248 ^ x216 ;
  assign n7601 = n7031 & n7032 ;
  assign n7606 = n7602 ^ n7601 ;
  assign n7627 = n7613 ^ n7606 ;
  assign n7708 = n7659 ^ n7627 ;
  assign n7029 = x119 ^ x87 ;
  assign n7030 = x247 ^ x215 ;
  assign n7522 = n7029 & n7030 ;
  assign n7027 = x118 ^ x86 ;
  assign n7028 = x246 ^ x214 ;
  assign n7521 = n7027 & n7028 ;
  assign n7526 = n7522 ^ n7521 ;
  assign n7025 = x117 ^ x85 ;
  assign n7026 = x245 ^ x213 ;
  assign n7515 = n7025 & n7026 ;
  assign n7023 = x116 ^ x84 ;
  assign n7024 = x244 ^ x212 ;
  assign n7514 = n7023 & n7024 ;
  assign n7519 = n7515 ^ n7514 ;
  assign n7540 = n7526 ^ n7519 ;
  assign n7021 = x115 ^ x83 ;
  assign n7022 = x243 ^ x211 ;
  assign n7490 = n7021 & n7022 ;
  assign n7019 = x114 ^ x82 ;
  assign n7020 = x242 ^ x210 ;
  assign n7489 = n7019 & n7020 ;
  assign n7494 = n7490 ^ n7489 ;
  assign n7017 = x113 ^ x81 ;
  assign n7018 = x241 ^ x209 ;
  assign n7483 = n7017 & n7018 ;
  assign n7015 = x112 ^ x80 ;
  assign n7016 = x240 ^ x208 ;
  assign n7482 = n7015 & n7016 ;
  assign n7487 = n7483 ^ n7482 ;
  assign n7508 = n7494 ^ n7487 ;
  assign n7589 = n7540 ^ n7508 ;
  assign n7862 = n7708 ^ n7589 ;
  assign n7013 = x111 ^ x79 ;
  assign n7014 = x239 ^ x207 ;
  assign n7237 = n7013 & n7014 ;
  assign n7011 = x110 ^ x78 ;
  assign n7012 = x238 ^ x206 ;
  assign n7236 = n7011 & n7012 ;
  assign n7241 = n7237 ^ n7236 ;
  assign n7009 = x109 ^ x77 ;
  assign n7010 = x237 ^ x205 ;
  assign n7230 = n7009 & n7010 ;
  assign n7007 = x108 ^ x76 ;
  assign n7008 = x236 ^ x204 ;
  assign n7229 = n7007 & n7008 ;
  assign n7234 = n7230 ^ n7229 ;
  assign n7255 = n7241 ^ n7234 ;
  assign n7005 = x107 ^ x75 ;
  assign n7006 = x235 ^ x203 ;
  assign n7205 = n7005 & n7006 ;
  assign n7003 = x106 ^ x74 ;
  assign n7004 = x234 ^ x202 ;
  assign n7204 = n7003 & n7004 ;
  assign n7209 = n7205 ^ n7204 ;
  assign n7001 = x105 ^ x73 ;
  assign n7002 = x233 ^ x201 ;
  assign n7198 = n7001 & n7002 ;
  assign n6999 = x104 ^ x72 ;
  assign n7000 = x232 ^ x200 ;
  assign n7197 = n6999 & n7000 ;
  assign n7202 = n7198 ^ n7197 ;
  assign n7223 = n7209 ^ n7202 ;
  assign n7304 = n7255 ^ n7223 ;
  assign n6997 = x103 ^ x71 ;
  assign n6998 = x231 ^ x199 ;
  assign n7118 = n6997 & n6998 ;
  assign n6995 = x102 ^ x70 ;
  assign n6996 = x230 ^ x198 ;
  assign n7117 = n6995 & n6996 ;
  assign n7122 = n7118 ^ n7117 ;
  assign n6993 = x101 ^ x69 ;
  assign n6994 = x229 ^ x197 ;
  assign n7111 = n6993 & n6994 ;
  assign n6991 = x100 ^ x68 ;
  assign n6992 = x228 ^ x196 ;
  assign n7110 = n6991 & n6992 ;
  assign n7115 = n7111 ^ n7110 ;
  assign n7136 = n7122 ^ n7115 ;
  assign n6989 = x99 ^ x67 ;
  assign n6990 = x227 ^ x195 ;
  assign n7086 = n6989 & n6990 ;
  assign n6987 = x98 ^ x66 ;
  assign n6988 = x226 ^ x194 ;
  assign n7085 = n6987 & n6988 ;
  assign n7090 = n7086 ^ n7085 ;
  assign n6985 = x97 ^ x65 ;
  assign n6986 = x225 ^ x193 ;
  assign n7079 = n6985 & n6986 ;
  assign n6983 = x96 ^ x64 ;
  assign n6984 = x224 ^ x192 ;
  assign n7078 = n6983 & n6984 ;
  assign n7083 = n7079 ^ n7078 ;
  assign n7104 = n7090 ^ n7083 ;
  assign n7185 = n7136 ^ n7104 ;
  assign n7458 = n7304 ^ n7185 ;
  assign n8337 = n7862 ^ n7458 ;
  assign n8417 = n8385 ^ n8337 ;
  assign n8418 = n8417 ^ n6952 ;
  assign n2933 = x63 ^ x31 ;
  assign n2934 = x191 ^ x159 ;
  assign n3529 = n2933 & n2934 ;
  assign n2931 = x62 ^ x30 ;
  assign n2932 = x190 ^ x158 ;
  assign n3528 = n2931 & n2932 ;
  assign n3533 = n3529 ^ n3528 ;
  assign n2929 = x61 ^ x29 ;
  assign n2930 = x189 ^ x157 ;
  assign n3522 = n2929 & n2930 ;
  assign n2927 = x60 ^ x28 ;
  assign n2928 = x188 ^ x156 ;
  assign n3521 = n2927 & n2928 ;
  assign n3526 = n3522 ^ n3521 ;
  assign n3547 = n3533 ^ n3526 ;
  assign n2925 = x59 ^ x27 ;
  assign n2926 = x187 ^ x155 ;
  assign n3497 = n2925 & n2926 ;
  assign n2923 = x58 ^ x26 ;
  assign n2924 = x186 ^ x154 ;
  assign n3496 = n2923 & n2924 ;
  assign n3501 = n3497 ^ n3496 ;
  assign n2921 = x57 ^ x25 ;
  assign n2922 = x185 ^ x153 ;
  assign n3490 = n2921 & n2922 ;
  assign n2919 = x56 ^ x24 ;
  assign n2920 = x184 ^ x152 ;
  assign n3489 = n2919 & n2920 ;
  assign n3494 = n3490 ^ n3489 ;
  assign n3515 = n3501 ^ n3494 ;
  assign n3596 = n3547 ^ n3515 ;
  assign n2917 = x55 ^ x23 ;
  assign n2918 = x183 ^ x151 ;
  assign n3410 = n2917 & n2918 ;
  assign n2915 = x54 ^ x22 ;
  assign n2916 = x182 ^ x150 ;
  assign n3409 = n2915 & n2916 ;
  assign n3414 = n3410 ^ n3409 ;
  assign n2913 = x53 ^ x21 ;
  assign n2914 = x181 ^ x149 ;
  assign n3403 = n2913 & n2914 ;
  assign n2911 = x52 ^ x20 ;
  assign n2912 = x180 ^ x148 ;
  assign n3402 = n2911 & n2912 ;
  assign n3407 = n3403 ^ n3402 ;
  assign n3428 = n3414 ^ n3407 ;
  assign n2909 = x51 ^ x19 ;
  assign n2910 = x179 ^ x147 ;
  assign n3378 = n2909 & n2910 ;
  assign n2907 = x50 ^ x18 ;
  assign n2908 = x178 ^ x146 ;
  assign n3377 = n2907 & n2908 ;
  assign n3382 = n3378 ^ n3377 ;
  assign n2905 = x49 ^ x17 ;
  assign n2906 = x177 ^ x145 ;
  assign n3371 = n2905 & n2906 ;
  assign n2903 = x48 ^ x16 ;
  assign n2904 = x176 ^ x144 ;
  assign n3370 = n2903 & n2904 ;
  assign n3375 = n3371 ^ n3370 ;
  assign n3396 = n3382 ^ n3375 ;
  assign n3477 = n3428 ^ n3396 ;
  assign n3750 = n3596 ^ n3477 ;
  assign n2901 = x47 ^ x15 ;
  assign n2902 = x175 ^ x143 ;
  assign n3125 = n2901 & n2902 ;
  assign n2899 = x46 ^ x14 ;
  assign n2900 = x174 ^ x142 ;
  assign n3124 = n2899 & n2900 ;
  assign n3129 = n3125 ^ n3124 ;
  assign n2897 = x45 ^ x13 ;
  assign n2898 = x173 ^ x141 ;
  assign n3118 = n2897 & n2898 ;
  assign n2895 = x44 ^ x12 ;
  assign n2896 = x172 ^ x140 ;
  assign n3117 = n2895 & n2896 ;
  assign n3122 = n3118 ^ n3117 ;
  assign n3143 = n3129 ^ n3122 ;
  assign n2893 = x43 ^ x11 ;
  assign n2894 = x171 ^ x139 ;
  assign n3093 = n2893 & n2894 ;
  assign n2891 = x42 ^ x10 ;
  assign n2892 = x170 ^ x138 ;
  assign n3092 = n2891 & n2892 ;
  assign n3097 = n3093 ^ n3092 ;
  assign n2889 = x41 ^ x9 ;
  assign n2890 = x169 ^ x137 ;
  assign n3086 = n2889 & n2890 ;
  assign n2887 = x40 ^ x8 ;
  assign n2888 = x168 ^ x136 ;
  assign n3085 = n2887 & n2888 ;
  assign n3090 = n3086 ^ n3085 ;
  assign n3111 = n3097 ^ n3090 ;
  assign n3192 = n3143 ^ n3111 ;
  assign n2885 = x39 ^ x7 ;
  assign n2886 = x167 ^ x135 ;
  assign n3006 = n2885 & n2886 ;
  assign n2883 = x38 ^ x6 ;
  assign n2884 = x166 ^ x134 ;
  assign n3005 = n2883 & n2884 ;
  assign n3010 = n3006 ^ n3005 ;
  assign n2881 = x37 ^ x5 ;
  assign n2882 = x165 ^ x133 ;
  assign n2999 = n2881 & n2882 ;
  assign n2879 = x36 ^ x4 ;
  assign n2880 = x164 ^ x132 ;
  assign n2998 = n2879 & n2880 ;
  assign n3003 = n2999 ^ n2998 ;
  assign n3024 = n3010 ^ n3003 ;
  assign n2877 = x35 ^ x3 ;
  assign n2878 = x163 ^ x131 ;
  assign n2974 = n2877 & n2878 ;
  assign n2875 = x34 ^ x2 ;
  assign n2876 = x162 ^ x130 ;
  assign n2973 = n2875 & n2876 ;
  assign n2978 = n2974 ^ n2973 ;
  assign n2873 = x33 ^ x1 ;
  assign n2874 = x161 ^ x129 ;
  assign n2967 = n2873 & n2874 ;
  assign n2871 = x32 ^ x0 ;
  assign n2872 = x160 ^ x128 ;
  assign n2966 = n2871 & n2872 ;
  assign n2971 = n2967 ^ n2966 ;
  assign n2992 = n2978 ^ n2971 ;
  assign n3073 = n3024 ^ n2992 ;
  assign n3346 = n3192 ^ n3073 ;
  assign n4225 = n3750 ^ n3346 ;
  assign n4305 = n4273 ^ n4225 ;
  assign n4306 = n4305 ^ n2840 ;
  assign n12816 = n8418 ^ n4306 ;
  assign n7642 = n7045 ^ n7043 ;
  assign n7643 = n7046 ^ n7044 ;
  assign n7644 = n7642 & n7643 ;
  assign n7646 = n7644 ^ n7640 ;
  assign n7635 = n7041 ^ n7039 ;
  assign n7636 = n7042 ^ n7040 ;
  assign n7637 = n7635 & n7636 ;
  assign n7639 = n7637 ^ n7633 ;
  assign n7660 = n7646 ^ n7639 ;
  assign n7610 = n7037 ^ n7035 ;
  assign n7611 = n7038 ^ n7036 ;
  assign n7612 = n7610 & n7611 ;
  assign n7614 = n7612 ^ n7608 ;
  assign n7603 = n7033 ^ n7031 ;
  assign n7604 = n7034 ^ n7032 ;
  assign n7605 = n7603 & n7604 ;
  assign n7607 = n7605 ^ n7601 ;
  assign n7628 = n7614 ^ n7607 ;
  assign n7709 = n7660 ^ n7628 ;
  assign n7523 = n7029 ^ n7027 ;
  assign n7524 = n7030 ^ n7028 ;
  assign n7525 = n7523 & n7524 ;
  assign n7527 = n7525 ^ n7521 ;
  assign n7516 = n7025 ^ n7023 ;
  assign n7517 = n7026 ^ n7024 ;
  assign n7518 = n7516 & n7517 ;
  assign n7520 = n7518 ^ n7514 ;
  assign n7541 = n7527 ^ n7520 ;
  assign n7491 = n7021 ^ n7019 ;
  assign n7492 = n7022 ^ n7020 ;
  assign n7493 = n7491 & n7492 ;
  assign n7495 = n7493 ^ n7489 ;
  assign n7484 = n7017 ^ n7015 ;
  assign n7485 = n7018 ^ n7016 ;
  assign n7486 = n7484 & n7485 ;
  assign n7488 = n7486 ^ n7482 ;
  assign n7509 = n7495 ^ n7488 ;
  assign n7590 = n7541 ^ n7509 ;
  assign n7863 = n7709 ^ n7590 ;
  assign n7238 = n7013 ^ n7011 ;
  assign n7239 = n7014 ^ n7012 ;
  assign n7240 = n7238 & n7239 ;
  assign n7242 = n7240 ^ n7236 ;
  assign n7231 = n7009 ^ n7007 ;
  assign n7232 = n7010 ^ n7008 ;
  assign n7233 = n7231 & n7232 ;
  assign n7235 = n7233 ^ n7229 ;
  assign n7256 = n7242 ^ n7235 ;
  assign n7206 = n7005 ^ n7003 ;
  assign n7207 = n7006 ^ n7004 ;
  assign n7208 = n7206 & n7207 ;
  assign n7210 = n7208 ^ n7204 ;
  assign n7199 = n7001 ^ n6999 ;
  assign n7200 = n7002 ^ n7000 ;
  assign n7201 = n7199 & n7200 ;
  assign n7203 = n7201 ^ n7197 ;
  assign n7224 = n7210 ^ n7203 ;
  assign n7305 = n7256 ^ n7224 ;
  assign n7119 = n6997 ^ n6995 ;
  assign n7120 = n6998 ^ n6996 ;
  assign n7121 = n7119 & n7120 ;
  assign n7123 = n7121 ^ n7117 ;
  assign n7112 = n6993 ^ n6991 ;
  assign n7113 = n6994 ^ n6992 ;
  assign n7114 = n7112 & n7113 ;
  assign n7116 = n7114 ^ n7110 ;
  assign n7137 = n7123 ^ n7116 ;
  assign n7087 = n6989 ^ n6987 ;
  assign n7088 = n6990 ^ n6988 ;
  assign n7089 = n7087 & n7088 ;
  assign n7091 = n7089 ^ n7085 ;
  assign n7080 = n6985 ^ n6983 ;
  assign n7081 = n6986 ^ n6984 ;
  assign n7082 = n7080 & n7081 ;
  assign n7084 = n7082 ^ n7078 ;
  assign n7105 = n7091 ^ n7084 ;
  assign n7186 = n7137 ^ n7105 ;
  assign n7459 = n7305 ^ n7186 ;
  assign n8338 = n7863 ^ n7459 ;
  assign n8419 = n8386 ^ n8338 ;
  assign n8420 = n8419 ^ n6954 ;
  assign n3530 = n2933 ^ n2931 ;
  assign n3531 = n2934 ^ n2932 ;
  assign n3532 = n3530 & n3531 ;
  assign n3534 = n3532 ^ n3528 ;
  assign n3523 = n2929 ^ n2927 ;
  assign n3524 = n2930 ^ n2928 ;
  assign n3525 = n3523 & n3524 ;
  assign n3527 = n3525 ^ n3521 ;
  assign n3548 = n3534 ^ n3527 ;
  assign n3498 = n2925 ^ n2923 ;
  assign n3499 = n2926 ^ n2924 ;
  assign n3500 = n3498 & n3499 ;
  assign n3502 = n3500 ^ n3496 ;
  assign n3491 = n2921 ^ n2919 ;
  assign n3492 = n2922 ^ n2920 ;
  assign n3493 = n3491 & n3492 ;
  assign n3495 = n3493 ^ n3489 ;
  assign n3516 = n3502 ^ n3495 ;
  assign n3597 = n3548 ^ n3516 ;
  assign n3411 = n2917 ^ n2915 ;
  assign n3412 = n2918 ^ n2916 ;
  assign n3413 = n3411 & n3412 ;
  assign n3415 = n3413 ^ n3409 ;
  assign n3404 = n2913 ^ n2911 ;
  assign n3405 = n2914 ^ n2912 ;
  assign n3406 = n3404 & n3405 ;
  assign n3408 = n3406 ^ n3402 ;
  assign n3429 = n3415 ^ n3408 ;
  assign n3379 = n2909 ^ n2907 ;
  assign n3380 = n2910 ^ n2908 ;
  assign n3381 = n3379 & n3380 ;
  assign n3383 = n3381 ^ n3377 ;
  assign n3372 = n2905 ^ n2903 ;
  assign n3373 = n2906 ^ n2904 ;
  assign n3374 = n3372 & n3373 ;
  assign n3376 = n3374 ^ n3370 ;
  assign n3397 = n3383 ^ n3376 ;
  assign n3478 = n3429 ^ n3397 ;
  assign n3751 = n3597 ^ n3478 ;
  assign n3126 = n2901 ^ n2899 ;
  assign n3127 = n2902 ^ n2900 ;
  assign n3128 = n3126 & n3127 ;
  assign n3130 = n3128 ^ n3124 ;
  assign n3119 = n2897 ^ n2895 ;
  assign n3120 = n2898 ^ n2896 ;
  assign n3121 = n3119 & n3120 ;
  assign n3123 = n3121 ^ n3117 ;
  assign n3144 = n3130 ^ n3123 ;
  assign n3094 = n2893 ^ n2891 ;
  assign n3095 = n2894 ^ n2892 ;
  assign n3096 = n3094 & n3095 ;
  assign n3098 = n3096 ^ n3092 ;
  assign n3087 = n2889 ^ n2887 ;
  assign n3088 = n2890 ^ n2888 ;
  assign n3089 = n3087 & n3088 ;
  assign n3091 = n3089 ^ n3085 ;
  assign n3112 = n3098 ^ n3091 ;
  assign n3193 = n3144 ^ n3112 ;
  assign n3007 = n2885 ^ n2883 ;
  assign n3008 = n2886 ^ n2884 ;
  assign n3009 = n3007 & n3008 ;
  assign n3011 = n3009 ^ n3005 ;
  assign n3000 = n2881 ^ n2879 ;
  assign n3001 = n2882 ^ n2880 ;
  assign n3002 = n3000 & n3001 ;
  assign n3004 = n3002 ^ n2998 ;
  assign n3025 = n3011 ^ n3004 ;
  assign n2975 = n2877 ^ n2875 ;
  assign n2976 = n2878 ^ n2876 ;
  assign n2977 = n2975 & n2976 ;
  assign n2979 = n2977 ^ n2973 ;
  assign n2968 = n2873 ^ n2871 ;
  assign n2969 = n2874 ^ n2872 ;
  assign n2970 = n2968 & n2969 ;
  assign n2972 = n2970 ^ n2966 ;
  assign n2993 = n2979 ^ n2972 ;
  assign n3074 = n3025 ^ n2993 ;
  assign n3347 = n3193 ^ n3074 ;
  assign n4226 = n3751 ^ n3347 ;
  assign n4307 = n4274 ^ n4226 ;
  assign n4308 = n4307 ^ n2842 ;
  assign n12817 = n8420 ^ n4308 ;
  assign n7649 = n7045 ^ n7041 ;
  assign n7650 = n7046 ^ n7042 ;
  assign n7653 = n7649 & n7650 ;
  assign n7647 = n7043 ^ n7039 ;
  assign n7648 = n7044 ^ n7040 ;
  assign n7652 = n7647 & n7648 ;
  assign n7657 = n7653 ^ n7652 ;
  assign n7661 = n7659 ^ n7657 ;
  assign n7662 = n7661 ^ n7646 ;
  assign n7617 = n7037 ^ n7033 ;
  assign n7618 = n7038 ^ n7034 ;
  assign n7621 = n7617 & n7618 ;
  assign n7615 = n7035 ^ n7031 ;
  assign n7616 = n7036 ^ n7032 ;
  assign n7620 = n7615 & n7616 ;
  assign n7625 = n7621 ^ n7620 ;
  assign n7629 = n7627 ^ n7625 ;
  assign n7630 = n7629 ^ n7614 ;
  assign n7710 = n7662 ^ n7630 ;
  assign n7530 = n7029 ^ n7025 ;
  assign n7531 = n7030 ^ n7026 ;
  assign n7534 = n7530 & n7531 ;
  assign n7528 = n7027 ^ n7023 ;
  assign n7529 = n7028 ^ n7024 ;
  assign n7533 = n7528 & n7529 ;
  assign n7538 = n7534 ^ n7533 ;
  assign n7542 = n7540 ^ n7538 ;
  assign n7543 = n7542 ^ n7527 ;
  assign n7498 = n7021 ^ n7017 ;
  assign n7499 = n7022 ^ n7018 ;
  assign n7502 = n7498 & n7499 ;
  assign n7496 = n7019 ^ n7015 ;
  assign n7497 = n7020 ^ n7016 ;
  assign n7501 = n7496 & n7497 ;
  assign n7506 = n7502 ^ n7501 ;
  assign n7510 = n7508 ^ n7506 ;
  assign n7511 = n7510 ^ n7495 ;
  assign n7591 = n7543 ^ n7511 ;
  assign n7864 = n7710 ^ n7591 ;
  assign n7245 = n7013 ^ n7009 ;
  assign n7246 = n7014 ^ n7010 ;
  assign n7249 = n7245 & n7246 ;
  assign n7243 = n7011 ^ n7007 ;
  assign n7244 = n7012 ^ n7008 ;
  assign n7248 = n7243 & n7244 ;
  assign n7253 = n7249 ^ n7248 ;
  assign n7257 = n7255 ^ n7253 ;
  assign n7258 = n7257 ^ n7242 ;
  assign n7213 = n7005 ^ n7001 ;
  assign n7214 = n7006 ^ n7002 ;
  assign n7217 = n7213 & n7214 ;
  assign n7211 = n7003 ^ n6999 ;
  assign n7212 = n7004 ^ n7000 ;
  assign n7216 = n7211 & n7212 ;
  assign n7221 = n7217 ^ n7216 ;
  assign n7225 = n7223 ^ n7221 ;
  assign n7226 = n7225 ^ n7210 ;
  assign n7306 = n7258 ^ n7226 ;
  assign n7126 = n6997 ^ n6993 ;
  assign n7127 = n6998 ^ n6994 ;
  assign n7130 = n7126 & n7127 ;
  assign n7124 = n6995 ^ n6991 ;
  assign n7125 = n6996 ^ n6992 ;
  assign n7129 = n7124 & n7125 ;
  assign n7134 = n7130 ^ n7129 ;
  assign n7138 = n7136 ^ n7134 ;
  assign n7139 = n7138 ^ n7123 ;
  assign n7094 = n6989 ^ n6985 ;
  assign n7095 = n6990 ^ n6986 ;
  assign n7098 = n7094 & n7095 ;
  assign n7092 = n6987 ^ n6983 ;
  assign n7093 = n6988 ^ n6984 ;
  assign n7097 = n7092 & n7093 ;
  assign n7102 = n7098 ^ n7097 ;
  assign n7106 = n7104 ^ n7102 ;
  assign n7107 = n7106 ^ n7091 ;
  assign n7187 = n7139 ^ n7107 ;
  assign n7460 = n7306 ^ n7187 ;
  assign n8339 = n7864 ^ n7460 ;
  assign n8421 = n8387 ^ n8339 ;
  assign n8422 = n8421 ^ n6956 ;
  assign n3537 = n2933 ^ n2929 ;
  assign n3538 = n2934 ^ n2930 ;
  assign n3541 = n3537 & n3538 ;
  assign n3535 = n2931 ^ n2927 ;
  assign n3536 = n2932 ^ n2928 ;
  assign n3540 = n3535 & n3536 ;
  assign n3545 = n3541 ^ n3540 ;
  assign n3549 = n3547 ^ n3545 ;
  assign n3550 = n3549 ^ n3534 ;
  assign n3505 = n2925 ^ n2921 ;
  assign n3506 = n2926 ^ n2922 ;
  assign n3509 = n3505 & n3506 ;
  assign n3503 = n2923 ^ n2919 ;
  assign n3504 = n2924 ^ n2920 ;
  assign n3508 = n3503 & n3504 ;
  assign n3513 = n3509 ^ n3508 ;
  assign n3517 = n3515 ^ n3513 ;
  assign n3518 = n3517 ^ n3502 ;
  assign n3598 = n3550 ^ n3518 ;
  assign n3418 = n2917 ^ n2913 ;
  assign n3419 = n2918 ^ n2914 ;
  assign n3422 = n3418 & n3419 ;
  assign n3416 = n2915 ^ n2911 ;
  assign n3417 = n2916 ^ n2912 ;
  assign n3421 = n3416 & n3417 ;
  assign n3426 = n3422 ^ n3421 ;
  assign n3430 = n3428 ^ n3426 ;
  assign n3431 = n3430 ^ n3415 ;
  assign n3386 = n2909 ^ n2905 ;
  assign n3387 = n2910 ^ n2906 ;
  assign n3390 = n3386 & n3387 ;
  assign n3384 = n2907 ^ n2903 ;
  assign n3385 = n2908 ^ n2904 ;
  assign n3389 = n3384 & n3385 ;
  assign n3394 = n3390 ^ n3389 ;
  assign n3398 = n3396 ^ n3394 ;
  assign n3399 = n3398 ^ n3383 ;
  assign n3479 = n3431 ^ n3399 ;
  assign n3752 = n3598 ^ n3479 ;
  assign n3133 = n2901 ^ n2897 ;
  assign n3134 = n2902 ^ n2898 ;
  assign n3137 = n3133 & n3134 ;
  assign n3131 = n2899 ^ n2895 ;
  assign n3132 = n2900 ^ n2896 ;
  assign n3136 = n3131 & n3132 ;
  assign n3141 = n3137 ^ n3136 ;
  assign n3145 = n3143 ^ n3141 ;
  assign n3146 = n3145 ^ n3130 ;
  assign n3101 = n2893 ^ n2889 ;
  assign n3102 = n2894 ^ n2890 ;
  assign n3105 = n3101 & n3102 ;
  assign n3099 = n2891 ^ n2887 ;
  assign n3100 = n2892 ^ n2888 ;
  assign n3104 = n3099 & n3100 ;
  assign n3109 = n3105 ^ n3104 ;
  assign n3113 = n3111 ^ n3109 ;
  assign n3114 = n3113 ^ n3098 ;
  assign n3194 = n3146 ^ n3114 ;
  assign n3014 = n2885 ^ n2881 ;
  assign n3015 = n2886 ^ n2882 ;
  assign n3018 = n3014 & n3015 ;
  assign n3012 = n2883 ^ n2879 ;
  assign n3013 = n2884 ^ n2880 ;
  assign n3017 = n3012 & n3013 ;
  assign n3022 = n3018 ^ n3017 ;
  assign n3026 = n3024 ^ n3022 ;
  assign n3027 = n3026 ^ n3011 ;
  assign n2982 = n2877 ^ n2873 ;
  assign n2983 = n2878 ^ n2874 ;
  assign n2986 = n2982 & n2983 ;
  assign n2980 = n2875 ^ n2871 ;
  assign n2981 = n2876 ^ n2872 ;
  assign n2985 = n2980 & n2981 ;
  assign n2990 = n2986 ^ n2985 ;
  assign n2994 = n2992 ^ n2990 ;
  assign n2995 = n2994 ^ n2979 ;
  assign n3075 = n3027 ^ n2995 ;
  assign n3348 = n3194 ^ n3075 ;
  assign n4227 = n3752 ^ n3348 ;
  assign n4309 = n4275 ^ n4227 ;
  assign n4310 = n4309 ^ n2844 ;
  assign n12818 = n8422 ^ n4310 ;
  assign n7654 = n7649 ^ n7647 ;
  assign n7655 = n7650 ^ n7648 ;
  assign n7656 = n7654 & n7655 ;
  assign n7658 = n7656 ^ n7652 ;
  assign n7663 = n7660 ^ n7658 ;
  assign n7651 = n7646 ^ n7645 ;
  assign n7664 = n7663 ^ n7651 ;
  assign n7622 = n7617 ^ n7615 ;
  assign n7623 = n7618 ^ n7616 ;
  assign n7624 = n7622 & n7623 ;
  assign n7626 = n7624 ^ n7620 ;
  assign n7631 = n7628 ^ n7626 ;
  assign n7619 = n7614 ^ n7613 ;
  assign n7632 = n7631 ^ n7619 ;
  assign n7711 = n7664 ^ n7632 ;
  assign n7535 = n7530 ^ n7528 ;
  assign n7536 = n7531 ^ n7529 ;
  assign n7537 = n7535 & n7536 ;
  assign n7539 = n7537 ^ n7533 ;
  assign n7544 = n7541 ^ n7539 ;
  assign n7532 = n7527 ^ n7526 ;
  assign n7545 = n7544 ^ n7532 ;
  assign n7503 = n7498 ^ n7496 ;
  assign n7504 = n7499 ^ n7497 ;
  assign n7505 = n7503 & n7504 ;
  assign n7507 = n7505 ^ n7501 ;
  assign n7512 = n7509 ^ n7507 ;
  assign n7500 = n7495 ^ n7494 ;
  assign n7513 = n7512 ^ n7500 ;
  assign n7592 = n7545 ^ n7513 ;
  assign n7865 = n7711 ^ n7592 ;
  assign n7250 = n7245 ^ n7243 ;
  assign n7251 = n7246 ^ n7244 ;
  assign n7252 = n7250 & n7251 ;
  assign n7254 = n7252 ^ n7248 ;
  assign n7259 = n7256 ^ n7254 ;
  assign n7247 = n7242 ^ n7241 ;
  assign n7260 = n7259 ^ n7247 ;
  assign n7218 = n7213 ^ n7211 ;
  assign n7219 = n7214 ^ n7212 ;
  assign n7220 = n7218 & n7219 ;
  assign n7222 = n7220 ^ n7216 ;
  assign n7227 = n7224 ^ n7222 ;
  assign n7215 = n7210 ^ n7209 ;
  assign n7228 = n7227 ^ n7215 ;
  assign n7307 = n7260 ^ n7228 ;
  assign n7131 = n7126 ^ n7124 ;
  assign n7132 = n7127 ^ n7125 ;
  assign n7133 = n7131 & n7132 ;
  assign n7135 = n7133 ^ n7129 ;
  assign n7140 = n7137 ^ n7135 ;
  assign n7128 = n7123 ^ n7122 ;
  assign n7141 = n7140 ^ n7128 ;
  assign n7099 = n7094 ^ n7092 ;
  assign n7100 = n7095 ^ n7093 ;
  assign n7101 = n7099 & n7100 ;
  assign n7103 = n7101 ^ n7097 ;
  assign n7108 = n7105 ^ n7103 ;
  assign n7096 = n7091 ^ n7090 ;
  assign n7109 = n7108 ^ n7096 ;
  assign n7188 = n7141 ^ n7109 ;
  assign n7461 = n7307 ^ n7188 ;
  assign n8340 = n7865 ^ n7461 ;
  assign n8423 = n8388 ^ n8340 ;
  assign n8424 = n8423 ^ n6958 ;
  assign n3542 = n3537 ^ n3535 ;
  assign n3543 = n3538 ^ n3536 ;
  assign n3544 = n3542 & n3543 ;
  assign n3546 = n3544 ^ n3540 ;
  assign n3551 = n3548 ^ n3546 ;
  assign n3539 = n3534 ^ n3533 ;
  assign n3552 = n3551 ^ n3539 ;
  assign n3510 = n3505 ^ n3503 ;
  assign n3511 = n3506 ^ n3504 ;
  assign n3512 = n3510 & n3511 ;
  assign n3514 = n3512 ^ n3508 ;
  assign n3519 = n3516 ^ n3514 ;
  assign n3507 = n3502 ^ n3501 ;
  assign n3520 = n3519 ^ n3507 ;
  assign n3599 = n3552 ^ n3520 ;
  assign n3423 = n3418 ^ n3416 ;
  assign n3424 = n3419 ^ n3417 ;
  assign n3425 = n3423 & n3424 ;
  assign n3427 = n3425 ^ n3421 ;
  assign n3432 = n3429 ^ n3427 ;
  assign n3420 = n3415 ^ n3414 ;
  assign n3433 = n3432 ^ n3420 ;
  assign n3391 = n3386 ^ n3384 ;
  assign n3392 = n3387 ^ n3385 ;
  assign n3393 = n3391 & n3392 ;
  assign n3395 = n3393 ^ n3389 ;
  assign n3400 = n3397 ^ n3395 ;
  assign n3388 = n3383 ^ n3382 ;
  assign n3401 = n3400 ^ n3388 ;
  assign n3480 = n3433 ^ n3401 ;
  assign n3753 = n3599 ^ n3480 ;
  assign n3138 = n3133 ^ n3131 ;
  assign n3139 = n3134 ^ n3132 ;
  assign n3140 = n3138 & n3139 ;
  assign n3142 = n3140 ^ n3136 ;
  assign n3147 = n3144 ^ n3142 ;
  assign n3135 = n3130 ^ n3129 ;
  assign n3148 = n3147 ^ n3135 ;
  assign n3106 = n3101 ^ n3099 ;
  assign n3107 = n3102 ^ n3100 ;
  assign n3108 = n3106 & n3107 ;
  assign n3110 = n3108 ^ n3104 ;
  assign n3115 = n3112 ^ n3110 ;
  assign n3103 = n3098 ^ n3097 ;
  assign n3116 = n3115 ^ n3103 ;
  assign n3195 = n3148 ^ n3116 ;
  assign n3019 = n3014 ^ n3012 ;
  assign n3020 = n3015 ^ n3013 ;
  assign n3021 = n3019 & n3020 ;
  assign n3023 = n3021 ^ n3017 ;
  assign n3028 = n3025 ^ n3023 ;
  assign n3016 = n3011 ^ n3010 ;
  assign n3029 = n3028 ^ n3016 ;
  assign n2987 = n2982 ^ n2980 ;
  assign n2988 = n2983 ^ n2981 ;
  assign n2989 = n2987 & n2988 ;
  assign n2991 = n2989 ^ n2985 ;
  assign n2996 = n2993 ^ n2991 ;
  assign n2984 = n2979 ^ n2978 ;
  assign n2997 = n2996 ^ n2984 ;
  assign n3076 = n3029 ^ n2997 ;
  assign n3349 = n3195 ^ n3076 ;
  assign n4228 = n3753 ^ n3349 ;
  assign n4311 = n4276 ^ n4228 ;
  assign n4312 = n4311 ^ n2846 ;
  assign n12819 = n8424 ^ n4312 ;
  assign n7671 = n7045 ^ n7037 ;
  assign n7672 = n7046 ^ n7038 ;
  assign n7684 = n7671 & n7672 ;
  assign n7669 = n7043 ^ n7035 ;
  assign n7670 = n7044 ^ n7036 ;
  assign n7683 = n7669 & n7670 ;
  assign n7688 = n7684 ^ n7683 ;
  assign n7667 = n7041 ^ n7033 ;
  assign n7668 = n7042 ^ n7034 ;
  assign n7677 = n7667 & n7668 ;
  assign n7665 = n7039 ^ n7031 ;
  assign n7666 = n7040 ^ n7032 ;
  assign n7676 = n7665 & n7666 ;
  assign n7681 = n7677 ^ n7676 ;
  assign n7702 = n7688 ^ n7681 ;
  assign n7712 = n7708 ^ n7702 ;
  assign n7713 = n7712 ^ n7662 ;
  assign n7552 = n7029 ^ n7021 ;
  assign n7553 = n7030 ^ n7022 ;
  assign n7565 = n7552 & n7553 ;
  assign n7550 = n7027 ^ n7019 ;
  assign n7551 = n7028 ^ n7020 ;
  assign n7564 = n7550 & n7551 ;
  assign n7569 = n7565 ^ n7564 ;
  assign n7548 = n7025 ^ n7017 ;
  assign n7549 = n7026 ^ n7018 ;
  assign n7558 = n7548 & n7549 ;
  assign n7546 = n7023 ^ n7015 ;
  assign n7547 = n7024 ^ n7016 ;
  assign n7557 = n7546 & n7547 ;
  assign n7562 = n7558 ^ n7557 ;
  assign n7583 = n7569 ^ n7562 ;
  assign n7593 = n7589 ^ n7583 ;
  assign n7594 = n7593 ^ n7543 ;
  assign n7866 = n7713 ^ n7594 ;
  assign n7267 = n7013 ^ n7005 ;
  assign n7268 = n7014 ^ n7006 ;
  assign n7280 = n7267 & n7268 ;
  assign n7265 = n7011 ^ n7003 ;
  assign n7266 = n7012 ^ n7004 ;
  assign n7279 = n7265 & n7266 ;
  assign n7284 = n7280 ^ n7279 ;
  assign n7263 = n7009 ^ n7001 ;
  assign n7264 = n7010 ^ n7002 ;
  assign n7273 = n7263 & n7264 ;
  assign n7261 = n7007 ^ n6999 ;
  assign n7262 = n7008 ^ n7000 ;
  assign n7272 = n7261 & n7262 ;
  assign n7277 = n7273 ^ n7272 ;
  assign n7298 = n7284 ^ n7277 ;
  assign n7308 = n7304 ^ n7298 ;
  assign n7309 = n7308 ^ n7258 ;
  assign n7148 = n6997 ^ n6989 ;
  assign n7149 = n6998 ^ n6990 ;
  assign n7161 = n7148 & n7149 ;
  assign n7146 = n6995 ^ n6987 ;
  assign n7147 = n6996 ^ n6988 ;
  assign n7160 = n7146 & n7147 ;
  assign n7165 = n7161 ^ n7160 ;
  assign n7144 = n6993 ^ n6985 ;
  assign n7145 = n6994 ^ n6986 ;
  assign n7154 = n7144 & n7145 ;
  assign n7142 = n6991 ^ n6983 ;
  assign n7143 = n6992 ^ n6984 ;
  assign n7153 = n7142 & n7143 ;
  assign n7158 = n7154 ^ n7153 ;
  assign n7179 = n7165 ^ n7158 ;
  assign n7189 = n7185 ^ n7179 ;
  assign n7190 = n7189 ^ n7139 ;
  assign n7462 = n7309 ^ n7190 ;
  assign n8341 = n7866 ^ n7462 ;
  assign n8425 = n8389 ^ n8341 ;
  assign n8426 = n8425 ^ n6960 ;
  assign n3559 = n2933 ^ n2925 ;
  assign n3560 = n2934 ^ n2926 ;
  assign n3572 = n3559 & n3560 ;
  assign n3557 = n2931 ^ n2923 ;
  assign n3558 = n2932 ^ n2924 ;
  assign n3571 = n3557 & n3558 ;
  assign n3576 = n3572 ^ n3571 ;
  assign n3555 = n2929 ^ n2921 ;
  assign n3556 = n2930 ^ n2922 ;
  assign n3565 = n3555 & n3556 ;
  assign n3553 = n2927 ^ n2919 ;
  assign n3554 = n2928 ^ n2920 ;
  assign n3564 = n3553 & n3554 ;
  assign n3569 = n3565 ^ n3564 ;
  assign n3590 = n3576 ^ n3569 ;
  assign n3600 = n3596 ^ n3590 ;
  assign n3601 = n3600 ^ n3550 ;
  assign n3440 = n2917 ^ n2909 ;
  assign n3441 = n2918 ^ n2910 ;
  assign n3453 = n3440 & n3441 ;
  assign n3438 = n2915 ^ n2907 ;
  assign n3439 = n2916 ^ n2908 ;
  assign n3452 = n3438 & n3439 ;
  assign n3457 = n3453 ^ n3452 ;
  assign n3436 = n2913 ^ n2905 ;
  assign n3437 = n2914 ^ n2906 ;
  assign n3446 = n3436 & n3437 ;
  assign n3434 = n2911 ^ n2903 ;
  assign n3435 = n2912 ^ n2904 ;
  assign n3445 = n3434 & n3435 ;
  assign n3450 = n3446 ^ n3445 ;
  assign n3471 = n3457 ^ n3450 ;
  assign n3481 = n3477 ^ n3471 ;
  assign n3482 = n3481 ^ n3431 ;
  assign n3754 = n3601 ^ n3482 ;
  assign n3155 = n2901 ^ n2893 ;
  assign n3156 = n2902 ^ n2894 ;
  assign n3168 = n3155 & n3156 ;
  assign n3153 = n2899 ^ n2891 ;
  assign n3154 = n2900 ^ n2892 ;
  assign n3167 = n3153 & n3154 ;
  assign n3172 = n3168 ^ n3167 ;
  assign n3151 = n2897 ^ n2889 ;
  assign n3152 = n2898 ^ n2890 ;
  assign n3161 = n3151 & n3152 ;
  assign n3149 = n2895 ^ n2887 ;
  assign n3150 = n2896 ^ n2888 ;
  assign n3160 = n3149 & n3150 ;
  assign n3165 = n3161 ^ n3160 ;
  assign n3186 = n3172 ^ n3165 ;
  assign n3196 = n3192 ^ n3186 ;
  assign n3197 = n3196 ^ n3146 ;
  assign n3036 = n2885 ^ n2877 ;
  assign n3037 = n2886 ^ n2878 ;
  assign n3049 = n3036 & n3037 ;
  assign n3034 = n2883 ^ n2875 ;
  assign n3035 = n2884 ^ n2876 ;
  assign n3048 = n3034 & n3035 ;
  assign n3053 = n3049 ^ n3048 ;
  assign n3032 = n2881 ^ n2873 ;
  assign n3033 = n2882 ^ n2874 ;
  assign n3042 = n3032 & n3033 ;
  assign n3030 = n2879 ^ n2871 ;
  assign n3031 = n2880 ^ n2872 ;
  assign n3041 = n3030 & n3031 ;
  assign n3046 = n3042 ^ n3041 ;
  assign n3067 = n3053 ^ n3046 ;
  assign n3077 = n3073 ^ n3067 ;
  assign n3078 = n3077 ^ n3027 ;
  assign n3350 = n3197 ^ n3078 ;
  assign n4229 = n3754 ^ n3350 ;
  assign n4313 = n4277 ^ n4229 ;
  assign n4314 = n4313 ^ n2848 ;
  assign n12820 = n8426 ^ n4314 ;
  assign n7685 = n7671 ^ n7669 ;
  assign n7686 = n7672 ^ n7670 ;
  assign n7687 = n7685 & n7686 ;
  assign n7689 = n7687 ^ n7683 ;
  assign n7678 = n7667 ^ n7665 ;
  assign n7679 = n7668 ^ n7666 ;
  assign n7680 = n7678 & n7679 ;
  assign n7682 = n7680 ^ n7676 ;
  assign n7703 = n7689 ^ n7682 ;
  assign n7714 = n7709 ^ n7703 ;
  assign n7715 = n7714 ^ n7664 ;
  assign n7566 = n7552 ^ n7550 ;
  assign n7567 = n7553 ^ n7551 ;
  assign n7568 = n7566 & n7567 ;
  assign n7570 = n7568 ^ n7564 ;
  assign n7559 = n7548 ^ n7546 ;
  assign n7560 = n7549 ^ n7547 ;
  assign n7561 = n7559 & n7560 ;
  assign n7563 = n7561 ^ n7557 ;
  assign n7584 = n7570 ^ n7563 ;
  assign n7595 = n7590 ^ n7584 ;
  assign n7596 = n7595 ^ n7545 ;
  assign n7867 = n7715 ^ n7596 ;
  assign n7281 = n7267 ^ n7265 ;
  assign n7282 = n7268 ^ n7266 ;
  assign n7283 = n7281 & n7282 ;
  assign n7285 = n7283 ^ n7279 ;
  assign n7274 = n7263 ^ n7261 ;
  assign n7275 = n7264 ^ n7262 ;
  assign n7276 = n7274 & n7275 ;
  assign n7278 = n7276 ^ n7272 ;
  assign n7299 = n7285 ^ n7278 ;
  assign n7310 = n7305 ^ n7299 ;
  assign n7311 = n7310 ^ n7260 ;
  assign n7162 = n7148 ^ n7146 ;
  assign n7163 = n7149 ^ n7147 ;
  assign n7164 = n7162 & n7163 ;
  assign n7166 = n7164 ^ n7160 ;
  assign n7155 = n7144 ^ n7142 ;
  assign n7156 = n7145 ^ n7143 ;
  assign n7157 = n7155 & n7156 ;
  assign n7159 = n7157 ^ n7153 ;
  assign n7180 = n7166 ^ n7159 ;
  assign n7191 = n7186 ^ n7180 ;
  assign n7192 = n7191 ^ n7141 ;
  assign n7463 = n7311 ^ n7192 ;
  assign n8342 = n7867 ^ n7463 ;
  assign n8427 = n8390 ^ n8342 ;
  assign n8428 = n8427 ^ n6962 ;
  assign n3573 = n3559 ^ n3557 ;
  assign n3574 = n3560 ^ n3558 ;
  assign n3575 = n3573 & n3574 ;
  assign n3577 = n3575 ^ n3571 ;
  assign n3566 = n3555 ^ n3553 ;
  assign n3567 = n3556 ^ n3554 ;
  assign n3568 = n3566 & n3567 ;
  assign n3570 = n3568 ^ n3564 ;
  assign n3591 = n3577 ^ n3570 ;
  assign n3602 = n3597 ^ n3591 ;
  assign n3603 = n3602 ^ n3552 ;
  assign n3454 = n3440 ^ n3438 ;
  assign n3455 = n3441 ^ n3439 ;
  assign n3456 = n3454 & n3455 ;
  assign n3458 = n3456 ^ n3452 ;
  assign n3447 = n3436 ^ n3434 ;
  assign n3448 = n3437 ^ n3435 ;
  assign n3449 = n3447 & n3448 ;
  assign n3451 = n3449 ^ n3445 ;
  assign n3472 = n3458 ^ n3451 ;
  assign n3483 = n3478 ^ n3472 ;
  assign n3484 = n3483 ^ n3433 ;
  assign n3755 = n3603 ^ n3484 ;
  assign n3169 = n3155 ^ n3153 ;
  assign n3170 = n3156 ^ n3154 ;
  assign n3171 = n3169 & n3170 ;
  assign n3173 = n3171 ^ n3167 ;
  assign n3162 = n3151 ^ n3149 ;
  assign n3163 = n3152 ^ n3150 ;
  assign n3164 = n3162 & n3163 ;
  assign n3166 = n3164 ^ n3160 ;
  assign n3187 = n3173 ^ n3166 ;
  assign n3198 = n3193 ^ n3187 ;
  assign n3199 = n3198 ^ n3148 ;
  assign n3050 = n3036 ^ n3034 ;
  assign n3051 = n3037 ^ n3035 ;
  assign n3052 = n3050 & n3051 ;
  assign n3054 = n3052 ^ n3048 ;
  assign n3043 = n3032 ^ n3030 ;
  assign n3044 = n3033 ^ n3031 ;
  assign n3045 = n3043 & n3044 ;
  assign n3047 = n3045 ^ n3041 ;
  assign n3068 = n3054 ^ n3047 ;
  assign n3079 = n3074 ^ n3068 ;
  assign n3080 = n3079 ^ n3029 ;
  assign n3351 = n3199 ^ n3080 ;
  assign n4230 = n3755 ^ n3351 ;
  assign n4315 = n4278 ^ n4230 ;
  assign n4316 = n4315 ^ n2850 ;
  assign n12821 = n8428 ^ n4316 ;
  assign n7692 = n7671 ^ n7667 ;
  assign n7693 = n7672 ^ n7668 ;
  assign n7696 = n7692 & n7693 ;
  assign n7690 = n7669 ^ n7665 ;
  assign n7691 = n7670 ^ n7666 ;
  assign n7695 = n7690 & n7691 ;
  assign n7700 = n7696 ^ n7695 ;
  assign n7704 = n7702 ^ n7700 ;
  assign n7705 = n7704 ^ n7689 ;
  assign n7716 = n7710 ^ n7705 ;
  assign n7674 = n7664 ^ n7659 ;
  assign n7717 = n7716 ^ n7674 ;
  assign n7573 = n7552 ^ n7548 ;
  assign n7574 = n7553 ^ n7549 ;
  assign n7577 = n7573 & n7574 ;
  assign n7571 = n7550 ^ n7546 ;
  assign n7572 = n7551 ^ n7547 ;
  assign n7576 = n7571 & n7572 ;
  assign n7581 = n7577 ^ n7576 ;
  assign n7585 = n7583 ^ n7581 ;
  assign n7586 = n7585 ^ n7570 ;
  assign n7597 = n7591 ^ n7586 ;
  assign n7555 = n7545 ^ n7540 ;
  assign n7598 = n7597 ^ n7555 ;
  assign n7868 = n7717 ^ n7598 ;
  assign n7288 = n7267 ^ n7263 ;
  assign n7289 = n7268 ^ n7264 ;
  assign n7292 = n7288 & n7289 ;
  assign n7286 = n7265 ^ n7261 ;
  assign n7287 = n7266 ^ n7262 ;
  assign n7291 = n7286 & n7287 ;
  assign n7296 = n7292 ^ n7291 ;
  assign n7300 = n7298 ^ n7296 ;
  assign n7301 = n7300 ^ n7285 ;
  assign n7312 = n7306 ^ n7301 ;
  assign n7270 = n7260 ^ n7255 ;
  assign n7313 = n7312 ^ n7270 ;
  assign n7169 = n7148 ^ n7144 ;
  assign n7170 = n7149 ^ n7145 ;
  assign n7173 = n7169 & n7170 ;
  assign n7167 = n7146 ^ n7142 ;
  assign n7168 = n7147 ^ n7143 ;
  assign n7172 = n7167 & n7168 ;
  assign n7177 = n7173 ^ n7172 ;
  assign n7181 = n7179 ^ n7177 ;
  assign n7182 = n7181 ^ n7166 ;
  assign n7193 = n7187 ^ n7182 ;
  assign n7151 = n7141 ^ n7136 ;
  assign n7194 = n7193 ^ n7151 ;
  assign n7464 = n7313 ^ n7194 ;
  assign n8343 = n7868 ^ n7464 ;
  assign n8429 = n8391 ^ n8343 ;
  assign n8430 = n8429 ^ n6964 ;
  assign n3580 = n3559 ^ n3555 ;
  assign n3581 = n3560 ^ n3556 ;
  assign n3584 = n3580 & n3581 ;
  assign n3578 = n3557 ^ n3553 ;
  assign n3579 = n3558 ^ n3554 ;
  assign n3583 = n3578 & n3579 ;
  assign n3588 = n3584 ^ n3583 ;
  assign n3592 = n3590 ^ n3588 ;
  assign n3593 = n3592 ^ n3577 ;
  assign n3604 = n3598 ^ n3593 ;
  assign n3562 = n3552 ^ n3547 ;
  assign n3605 = n3604 ^ n3562 ;
  assign n3461 = n3440 ^ n3436 ;
  assign n3462 = n3441 ^ n3437 ;
  assign n3465 = n3461 & n3462 ;
  assign n3459 = n3438 ^ n3434 ;
  assign n3460 = n3439 ^ n3435 ;
  assign n3464 = n3459 & n3460 ;
  assign n3469 = n3465 ^ n3464 ;
  assign n3473 = n3471 ^ n3469 ;
  assign n3474 = n3473 ^ n3458 ;
  assign n3485 = n3479 ^ n3474 ;
  assign n3443 = n3433 ^ n3428 ;
  assign n3486 = n3485 ^ n3443 ;
  assign n3756 = n3605 ^ n3486 ;
  assign n3176 = n3155 ^ n3151 ;
  assign n3177 = n3156 ^ n3152 ;
  assign n3180 = n3176 & n3177 ;
  assign n3174 = n3153 ^ n3149 ;
  assign n3175 = n3154 ^ n3150 ;
  assign n3179 = n3174 & n3175 ;
  assign n3184 = n3180 ^ n3179 ;
  assign n3188 = n3186 ^ n3184 ;
  assign n3189 = n3188 ^ n3173 ;
  assign n3200 = n3194 ^ n3189 ;
  assign n3158 = n3148 ^ n3143 ;
  assign n3201 = n3200 ^ n3158 ;
  assign n3057 = n3036 ^ n3032 ;
  assign n3058 = n3037 ^ n3033 ;
  assign n3061 = n3057 & n3058 ;
  assign n3055 = n3034 ^ n3030 ;
  assign n3056 = n3035 ^ n3031 ;
  assign n3060 = n3055 & n3056 ;
  assign n3065 = n3061 ^ n3060 ;
  assign n3069 = n3067 ^ n3065 ;
  assign n3070 = n3069 ^ n3054 ;
  assign n3081 = n3075 ^ n3070 ;
  assign n3039 = n3029 ^ n3024 ;
  assign n3082 = n3081 ^ n3039 ;
  assign n3352 = n3201 ^ n3082 ;
  assign n4231 = n3756 ^ n3352 ;
  assign n4317 = n4279 ^ n4231 ;
  assign n4318 = n4317 ^ n2852 ;
  assign n12822 = n8430 ^ n4318 ;
  assign n7697 = n7692 ^ n7690 ;
  assign n7698 = n7693 ^ n7691 ;
  assign n7699 = n7697 & n7698 ;
  assign n7701 = n7699 ^ n7695 ;
  assign n7706 = n7703 ^ n7701 ;
  assign n7694 = n7689 ^ n7688 ;
  assign n7707 = n7706 ^ n7694 ;
  assign n7718 = n7711 ^ n7707 ;
  assign n7673 = n7664 ^ n7662 ;
  assign n7675 = n7673 ^ n7660 ;
  assign n7719 = n7718 ^ n7675 ;
  assign n7578 = n7573 ^ n7571 ;
  assign n7579 = n7574 ^ n7572 ;
  assign n7580 = n7578 & n7579 ;
  assign n7582 = n7580 ^ n7576 ;
  assign n7587 = n7584 ^ n7582 ;
  assign n7575 = n7570 ^ n7569 ;
  assign n7588 = n7587 ^ n7575 ;
  assign n7599 = n7592 ^ n7588 ;
  assign n7554 = n7545 ^ n7543 ;
  assign n7556 = n7554 ^ n7541 ;
  assign n7600 = n7599 ^ n7556 ;
  assign n7869 = n7719 ^ n7600 ;
  assign n7293 = n7288 ^ n7286 ;
  assign n7294 = n7289 ^ n7287 ;
  assign n7295 = n7293 & n7294 ;
  assign n7297 = n7295 ^ n7291 ;
  assign n7302 = n7299 ^ n7297 ;
  assign n7290 = n7285 ^ n7284 ;
  assign n7303 = n7302 ^ n7290 ;
  assign n7314 = n7307 ^ n7303 ;
  assign n7269 = n7260 ^ n7258 ;
  assign n7271 = n7269 ^ n7256 ;
  assign n7315 = n7314 ^ n7271 ;
  assign n7174 = n7169 ^ n7167 ;
  assign n7175 = n7170 ^ n7168 ;
  assign n7176 = n7174 & n7175 ;
  assign n7178 = n7176 ^ n7172 ;
  assign n7183 = n7180 ^ n7178 ;
  assign n7171 = n7166 ^ n7165 ;
  assign n7184 = n7183 ^ n7171 ;
  assign n7195 = n7188 ^ n7184 ;
  assign n7150 = n7141 ^ n7139 ;
  assign n7152 = n7150 ^ n7137 ;
  assign n7196 = n7195 ^ n7152 ;
  assign n7465 = n7315 ^ n7196 ;
  assign n8344 = n7869 ^ n7465 ;
  assign n8431 = n8392 ^ n8344 ;
  assign n8432 = n8431 ^ n6966 ;
  assign n3585 = n3580 ^ n3578 ;
  assign n3586 = n3581 ^ n3579 ;
  assign n3587 = n3585 & n3586 ;
  assign n3589 = n3587 ^ n3583 ;
  assign n3594 = n3591 ^ n3589 ;
  assign n3582 = n3577 ^ n3576 ;
  assign n3595 = n3594 ^ n3582 ;
  assign n3606 = n3599 ^ n3595 ;
  assign n3561 = n3552 ^ n3550 ;
  assign n3563 = n3561 ^ n3548 ;
  assign n3607 = n3606 ^ n3563 ;
  assign n3466 = n3461 ^ n3459 ;
  assign n3467 = n3462 ^ n3460 ;
  assign n3468 = n3466 & n3467 ;
  assign n3470 = n3468 ^ n3464 ;
  assign n3475 = n3472 ^ n3470 ;
  assign n3463 = n3458 ^ n3457 ;
  assign n3476 = n3475 ^ n3463 ;
  assign n3487 = n3480 ^ n3476 ;
  assign n3442 = n3433 ^ n3431 ;
  assign n3444 = n3442 ^ n3429 ;
  assign n3488 = n3487 ^ n3444 ;
  assign n3757 = n3607 ^ n3488 ;
  assign n3181 = n3176 ^ n3174 ;
  assign n3182 = n3177 ^ n3175 ;
  assign n3183 = n3181 & n3182 ;
  assign n3185 = n3183 ^ n3179 ;
  assign n3190 = n3187 ^ n3185 ;
  assign n3178 = n3173 ^ n3172 ;
  assign n3191 = n3190 ^ n3178 ;
  assign n3202 = n3195 ^ n3191 ;
  assign n3157 = n3148 ^ n3146 ;
  assign n3159 = n3157 ^ n3144 ;
  assign n3203 = n3202 ^ n3159 ;
  assign n3062 = n3057 ^ n3055 ;
  assign n3063 = n3058 ^ n3056 ;
  assign n3064 = n3062 & n3063 ;
  assign n3066 = n3064 ^ n3060 ;
  assign n3071 = n3068 ^ n3066 ;
  assign n3059 = n3054 ^ n3053 ;
  assign n3072 = n3071 ^ n3059 ;
  assign n3083 = n3076 ^ n3072 ;
  assign n3038 = n3029 ^ n3027 ;
  assign n3040 = n3038 ^ n3025 ;
  assign n3084 = n3083 ^ n3040 ;
  assign n3353 = n3203 ^ n3084 ;
  assign n4232 = n3757 ^ n3353 ;
  assign n4319 = n4280 ^ n4232 ;
  assign n4320 = n4319 ^ n2854 ;
  assign n12823 = n8432 ^ n4320 ;
  assign n7734 = n7045 ^ n7029 ;
  assign n7735 = n7046 ^ n7030 ;
  assign n7783 = n7734 & n7735 ;
  assign n7732 = n7043 ^ n7027 ;
  assign n7733 = n7044 ^ n7028 ;
  assign n7782 = n7732 & n7733 ;
  assign n7787 = n7783 ^ n7782 ;
  assign n7730 = n7041 ^ n7025 ;
  assign n7731 = n7042 ^ n7026 ;
  assign n7776 = n7730 & n7731 ;
  assign n7728 = n7039 ^ n7023 ;
  assign n7729 = n7040 ^ n7024 ;
  assign n7775 = n7728 & n7729 ;
  assign n7780 = n7776 ^ n7775 ;
  assign n7801 = n7787 ^ n7780 ;
  assign n7726 = n7037 ^ n7021 ;
  assign n7727 = n7038 ^ n7022 ;
  assign n7751 = n7726 & n7727 ;
  assign n7724 = n7035 ^ n7019 ;
  assign n7725 = n7036 ^ n7020 ;
  assign n7750 = n7724 & n7725 ;
  assign n7755 = n7751 ^ n7750 ;
  assign n7722 = n7033 ^ n7017 ;
  assign n7723 = n7034 ^ n7018 ;
  assign n7744 = n7722 & n7723 ;
  assign n7720 = n7031 ^ n7015 ;
  assign n7721 = n7032 ^ n7016 ;
  assign n7743 = n7720 & n7721 ;
  assign n7748 = n7744 ^ n7743 ;
  assign n7769 = n7755 ^ n7748 ;
  assign n7850 = n7801 ^ n7769 ;
  assign n7870 = n7862 ^ n7850 ;
  assign n7871 = n7870 ^ n7713 ;
  assign n7330 = n7013 ^ n6997 ;
  assign n7331 = n7014 ^ n6998 ;
  assign n7379 = n7330 & n7331 ;
  assign n7328 = n7011 ^ n6995 ;
  assign n7329 = n7012 ^ n6996 ;
  assign n7378 = n7328 & n7329 ;
  assign n7383 = n7379 ^ n7378 ;
  assign n7326 = n7009 ^ n6993 ;
  assign n7327 = n7010 ^ n6994 ;
  assign n7372 = n7326 & n7327 ;
  assign n7324 = n7007 ^ n6991 ;
  assign n7325 = n7008 ^ n6992 ;
  assign n7371 = n7324 & n7325 ;
  assign n7376 = n7372 ^ n7371 ;
  assign n7397 = n7383 ^ n7376 ;
  assign n7322 = n7005 ^ n6989 ;
  assign n7323 = n7006 ^ n6990 ;
  assign n7347 = n7322 & n7323 ;
  assign n7320 = n7003 ^ n6987 ;
  assign n7321 = n7004 ^ n6988 ;
  assign n7346 = n7320 & n7321 ;
  assign n7351 = n7347 ^ n7346 ;
  assign n7318 = n7001 ^ n6985 ;
  assign n7319 = n7002 ^ n6986 ;
  assign n7340 = n7318 & n7319 ;
  assign n7316 = n6999 ^ n6983 ;
  assign n7317 = n7000 ^ n6984 ;
  assign n7339 = n7316 & n7317 ;
  assign n7344 = n7340 ^ n7339 ;
  assign n7365 = n7351 ^ n7344 ;
  assign n7446 = n7397 ^ n7365 ;
  assign n7466 = n7458 ^ n7446 ;
  assign n7467 = n7466 ^ n7309 ;
  assign n8345 = n7871 ^ n7467 ;
  assign n8433 = n8393 ^ n8345 ;
  assign n8434 = n8433 ^ n6968 ;
  assign n3622 = n2933 ^ n2917 ;
  assign n3623 = n2934 ^ n2918 ;
  assign n3671 = n3622 & n3623 ;
  assign n3620 = n2931 ^ n2915 ;
  assign n3621 = n2932 ^ n2916 ;
  assign n3670 = n3620 & n3621 ;
  assign n3675 = n3671 ^ n3670 ;
  assign n3618 = n2929 ^ n2913 ;
  assign n3619 = n2930 ^ n2914 ;
  assign n3664 = n3618 & n3619 ;
  assign n3616 = n2927 ^ n2911 ;
  assign n3617 = n2928 ^ n2912 ;
  assign n3663 = n3616 & n3617 ;
  assign n3668 = n3664 ^ n3663 ;
  assign n3689 = n3675 ^ n3668 ;
  assign n3614 = n2925 ^ n2909 ;
  assign n3615 = n2926 ^ n2910 ;
  assign n3639 = n3614 & n3615 ;
  assign n3612 = n2923 ^ n2907 ;
  assign n3613 = n2924 ^ n2908 ;
  assign n3638 = n3612 & n3613 ;
  assign n3643 = n3639 ^ n3638 ;
  assign n3610 = n2921 ^ n2905 ;
  assign n3611 = n2922 ^ n2906 ;
  assign n3632 = n3610 & n3611 ;
  assign n3608 = n2919 ^ n2903 ;
  assign n3609 = n2920 ^ n2904 ;
  assign n3631 = n3608 & n3609 ;
  assign n3636 = n3632 ^ n3631 ;
  assign n3657 = n3643 ^ n3636 ;
  assign n3738 = n3689 ^ n3657 ;
  assign n3758 = n3750 ^ n3738 ;
  assign n3759 = n3758 ^ n3601 ;
  assign n3218 = n2901 ^ n2885 ;
  assign n3219 = n2902 ^ n2886 ;
  assign n3267 = n3218 & n3219 ;
  assign n3216 = n2899 ^ n2883 ;
  assign n3217 = n2900 ^ n2884 ;
  assign n3266 = n3216 & n3217 ;
  assign n3271 = n3267 ^ n3266 ;
  assign n3214 = n2897 ^ n2881 ;
  assign n3215 = n2898 ^ n2882 ;
  assign n3260 = n3214 & n3215 ;
  assign n3212 = n2895 ^ n2879 ;
  assign n3213 = n2896 ^ n2880 ;
  assign n3259 = n3212 & n3213 ;
  assign n3264 = n3260 ^ n3259 ;
  assign n3285 = n3271 ^ n3264 ;
  assign n3210 = n2893 ^ n2877 ;
  assign n3211 = n2894 ^ n2878 ;
  assign n3235 = n3210 & n3211 ;
  assign n3208 = n2891 ^ n2875 ;
  assign n3209 = n2892 ^ n2876 ;
  assign n3234 = n3208 & n3209 ;
  assign n3239 = n3235 ^ n3234 ;
  assign n3206 = n2889 ^ n2873 ;
  assign n3207 = n2890 ^ n2874 ;
  assign n3228 = n3206 & n3207 ;
  assign n3204 = n2887 ^ n2871 ;
  assign n3205 = n2888 ^ n2872 ;
  assign n3227 = n3204 & n3205 ;
  assign n3232 = n3228 ^ n3227 ;
  assign n3253 = n3239 ^ n3232 ;
  assign n3334 = n3285 ^ n3253 ;
  assign n3354 = n3346 ^ n3334 ;
  assign n3355 = n3354 ^ n3197 ;
  assign n4233 = n3759 ^ n3355 ;
  assign n4321 = n4281 ^ n4233 ;
  assign n4322 = n4321 ^ n2856 ;
  assign n12824 = n8434 ^ n4322 ;
  assign n7784 = n7734 ^ n7732 ;
  assign n7785 = n7735 ^ n7733 ;
  assign n7786 = n7784 & n7785 ;
  assign n7788 = n7786 ^ n7782 ;
  assign n7777 = n7730 ^ n7728 ;
  assign n7778 = n7731 ^ n7729 ;
  assign n7779 = n7777 & n7778 ;
  assign n7781 = n7779 ^ n7775 ;
  assign n7802 = n7788 ^ n7781 ;
  assign n7752 = n7726 ^ n7724 ;
  assign n7753 = n7727 ^ n7725 ;
  assign n7754 = n7752 & n7753 ;
  assign n7756 = n7754 ^ n7750 ;
  assign n7745 = n7722 ^ n7720 ;
  assign n7746 = n7723 ^ n7721 ;
  assign n7747 = n7745 & n7746 ;
  assign n7749 = n7747 ^ n7743 ;
  assign n7770 = n7756 ^ n7749 ;
  assign n7851 = n7802 ^ n7770 ;
  assign n7872 = n7863 ^ n7851 ;
  assign n7873 = n7872 ^ n7715 ;
  assign n7380 = n7330 ^ n7328 ;
  assign n7381 = n7331 ^ n7329 ;
  assign n7382 = n7380 & n7381 ;
  assign n7384 = n7382 ^ n7378 ;
  assign n7373 = n7326 ^ n7324 ;
  assign n7374 = n7327 ^ n7325 ;
  assign n7375 = n7373 & n7374 ;
  assign n7377 = n7375 ^ n7371 ;
  assign n7398 = n7384 ^ n7377 ;
  assign n7348 = n7322 ^ n7320 ;
  assign n7349 = n7323 ^ n7321 ;
  assign n7350 = n7348 & n7349 ;
  assign n7352 = n7350 ^ n7346 ;
  assign n7341 = n7318 ^ n7316 ;
  assign n7342 = n7319 ^ n7317 ;
  assign n7343 = n7341 & n7342 ;
  assign n7345 = n7343 ^ n7339 ;
  assign n7366 = n7352 ^ n7345 ;
  assign n7447 = n7398 ^ n7366 ;
  assign n7468 = n7459 ^ n7447 ;
  assign n7469 = n7468 ^ n7311 ;
  assign n8346 = n7873 ^ n7469 ;
  assign n8435 = n8394 ^ n8346 ;
  assign n8436 = n8435 ^ n6970 ;
  assign n3672 = n3622 ^ n3620 ;
  assign n3673 = n3623 ^ n3621 ;
  assign n3674 = n3672 & n3673 ;
  assign n3676 = n3674 ^ n3670 ;
  assign n3665 = n3618 ^ n3616 ;
  assign n3666 = n3619 ^ n3617 ;
  assign n3667 = n3665 & n3666 ;
  assign n3669 = n3667 ^ n3663 ;
  assign n3690 = n3676 ^ n3669 ;
  assign n3640 = n3614 ^ n3612 ;
  assign n3641 = n3615 ^ n3613 ;
  assign n3642 = n3640 & n3641 ;
  assign n3644 = n3642 ^ n3638 ;
  assign n3633 = n3610 ^ n3608 ;
  assign n3634 = n3611 ^ n3609 ;
  assign n3635 = n3633 & n3634 ;
  assign n3637 = n3635 ^ n3631 ;
  assign n3658 = n3644 ^ n3637 ;
  assign n3739 = n3690 ^ n3658 ;
  assign n3760 = n3751 ^ n3739 ;
  assign n3761 = n3760 ^ n3603 ;
  assign n3268 = n3218 ^ n3216 ;
  assign n3269 = n3219 ^ n3217 ;
  assign n3270 = n3268 & n3269 ;
  assign n3272 = n3270 ^ n3266 ;
  assign n3261 = n3214 ^ n3212 ;
  assign n3262 = n3215 ^ n3213 ;
  assign n3263 = n3261 & n3262 ;
  assign n3265 = n3263 ^ n3259 ;
  assign n3286 = n3272 ^ n3265 ;
  assign n3236 = n3210 ^ n3208 ;
  assign n3237 = n3211 ^ n3209 ;
  assign n3238 = n3236 & n3237 ;
  assign n3240 = n3238 ^ n3234 ;
  assign n3229 = n3206 ^ n3204 ;
  assign n3230 = n3207 ^ n3205 ;
  assign n3231 = n3229 & n3230 ;
  assign n3233 = n3231 ^ n3227 ;
  assign n3254 = n3240 ^ n3233 ;
  assign n3335 = n3286 ^ n3254 ;
  assign n3356 = n3347 ^ n3335 ;
  assign n3357 = n3356 ^ n3199 ;
  assign n4234 = n3761 ^ n3357 ;
  assign n4323 = n4282 ^ n4234 ;
  assign n4324 = n4323 ^ n2858 ;
  assign n12825 = n8436 ^ n4324 ;
  assign n7791 = n7734 ^ n7730 ;
  assign n7792 = n7735 ^ n7731 ;
  assign n7795 = n7791 & n7792 ;
  assign n7789 = n7732 ^ n7728 ;
  assign n7790 = n7733 ^ n7729 ;
  assign n7794 = n7789 & n7790 ;
  assign n7799 = n7795 ^ n7794 ;
  assign n7803 = n7801 ^ n7799 ;
  assign n7804 = n7803 ^ n7788 ;
  assign n7759 = n7726 ^ n7722 ;
  assign n7760 = n7727 ^ n7723 ;
  assign n7763 = n7759 & n7760 ;
  assign n7757 = n7724 ^ n7720 ;
  assign n7758 = n7725 ^ n7721 ;
  assign n7762 = n7757 & n7758 ;
  assign n7767 = n7763 ^ n7762 ;
  assign n7771 = n7769 ^ n7767 ;
  assign n7772 = n7771 ^ n7756 ;
  assign n7852 = n7804 ^ n7772 ;
  assign n7874 = n7864 ^ n7852 ;
  assign n7875 = n7874 ^ n7717 ;
  assign n7387 = n7330 ^ n7326 ;
  assign n7388 = n7331 ^ n7327 ;
  assign n7391 = n7387 & n7388 ;
  assign n7385 = n7328 ^ n7324 ;
  assign n7386 = n7329 ^ n7325 ;
  assign n7390 = n7385 & n7386 ;
  assign n7395 = n7391 ^ n7390 ;
  assign n7399 = n7397 ^ n7395 ;
  assign n7400 = n7399 ^ n7384 ;
  assign n7355 = n7322 ^ n7318 ;
  assign n7356 = n7323 ^ n7319 ;
  assign n7359 = n7355 & n7356 ;
  assign n7353 = n7320 ^ n7316 ;
  assign n7354 = n7321 ^ n7317 ;
  assign n7358 = n7353 & n7354 ;
  assign n7363 = n7359 ^ n7358 ;
  assign n7367 = n7365 ^ n7363 ;
  assign n7368 = n7367 ^ n7352 ;
  assign n7448 = n7400 ^ n7368 ;
  assign n7470 = n7460 ^ n7448 ;
  assign n7471 = n7470 ^ n7313 ;
  assign n8347 = n7875 ^ n7471 ;
  assign n8437 = n8395 ^ n8347 ;
  assign n8438 = n8437 ^ n6972 ;
  assign n3679 = n3622 ^ n3618 ;
  assign n3680 = n3623 ^ n3619 ;
  assign n3683 = n3679 & n3680 ;
  assign n3677 = n3620 ^ n3616 ;
  assign n3678 = n3621 ^ n3617 ;
  assign n3682 = n3677 & n3678 ;
  assign n3687 = n3683 ^ n3682 ;
  assign n3691 = n3689 ^ n3687 ;
  assign n3692 = n3691 ^ n3676 ;
  assign n3647 = n3614 ^ n3610 ;
  assign n3648 = n3615 ^ n3611 ;
  assign n3651 = n3647 & n3648 ;
  assign n3645 = n3612 ^ n3608 ;
  assign n3646 = n3613 ^ n3609 ;
  assign n3650 = n3645 & n3646 ;
  assign n3655 = n3651 ^ n3650 ;
  assign n3659 = n3657 ^ n3655 ;
  assign n3660 = n3659 ^ n3644 ;
  assign n3740 = n3692 ^ n3660 ;
  assign n3762 = n3752 ^ n3740 ;
  assign n3763 = n3762 ^ n3605 ;
  assign n3275 = n3218 ^ n3214 ;
  assign n3276 = n3219 ^ n3215 ;
  assign n3279 = n3275 & n3276 ;
  assign n3273 = n3216 ^ n3212 ;
  assign n3274 = n3217 ^ n3213 ;
  assign n3278 = n3273 & n3274 ;
  assign n3283 = n3279 ^ n3278 ;
  assign n3287 = n3285 ^ n3283 ;
  assign n3288 = n3287 ^ n3272 ;
  assign n3243 = n3210 ^ n3206 ;
  assign n3244 = n3211 ^ n3207 ;
  assign n3247 = n3243 & n3244 ;
  assign n3241 = n3208 ^ n3204 ;
  assign n3242 = n3209 ^ n3205 ;
  assign n3246 = n3241 & n3242 ;
  assign n3251 = n3247 ^ n3246 ;
  assign n3255 = n3253 ^ n3251 ;
  assign n3256 = n3255 ^ n3240 ;
  assign n3336 = n3288 ^ n3256 ;
  assign n3358 = n3348 ^ n3336 ;
  assign n3359 = n3358 ^ n3201 ;
  assign n4235 = n3763 ^ n3359 ;
  assign n4325 = n4283 ^ n4235 ;
  assign n4326 = n4325 ^ n2860 ;
  assign n12826 = n8438 ^ n4326 ;
  assign n7796 = n7791 ^ n7789 ;
  assign n7797 = n7792 ^ n7790 ;
  assign n7798 = n7796 & n7797 ;
  assign n7800 = n7798 ^ n7794 ;
  assign n7805 = n7802 ^ n7800 ;
  assign n7793 = n7788 ^ n7787 ;
  assign n7806 = n7805 ^ n7793 ;
  assign n7764 = n7759 ^ n7757 ;
  assign n7765 = n7760 ^ n7758 ;
  assign n7766 = n7764 & n7765 ;
  assign n7768 = n7766 ^ n7762 ;
  assign n7773 = n7770 ^ n7768 ;
  assign n7761 = n7756 ^ n7755 ;
  assign n7774 = n7773 ^ n7761 ;
  assign n7853 = n7806 ^ n7774 ;
  assign n7876 = n7865 ^ n7853 ;
  assign n7877 = n7876 ^ n7719 ;
  assign n7392 = n7387 ^ n7385 ;
  assign n7393 = n7388 ^ n7386 ;
  assign n7394 = n7392 & n7393 ;
  assign n7396 = n7394 ^ n7390 ;
  assign n7401 = n7398 ^ n7396 ;
  assign n7389 = n7384 ^ n7383 ;
  assign n7402 = n7401 ^ n7389 ;
  assign n7360 = n7355 ^ n7353 ;
  assign n7361 = n7356 ^ n7354 ;
  assign n7362 = n7360 & n7361 ;
  assign n7364 = n7362 ^ n7358 ;
  assign n7369 = n7366 ^ n7364 ;
  assign n7357 = n7352 ^ n7351 ;
  assign n7370 = n7369 ^ n7357 ;
  assign n7449 = n7402 ^ n7370 ;
  assign n7472 = n7461 ^ n7449 ;
  assign n7473 = n7472 ^ n7315 ;
  assign n8348 = n7877 ^ n7473 ;
  assign n8439 = n8396 ^ n8348 ;
  assign n8440 = n8439 ^ n6974 ;
  assign n3684 = n3679 ^ n3677 ;
  assign n3685 = n3680 ^ n3678 ;
  assign n3686 = n3684 & n3685 ;
  assign n3688 = n3686 ^ n3682 ;
  assign n3693 = n3690 ^ n3688 ;
  assign n3681 = n3676 ^ n3675 ;
  assign n3694 = n3693 ^ n3681 ;
  assign n3652 = n3647 ^ n3645 ;
  assign n3653 = n3648 ^ n3646 ;
  assign n3654 = n3652 & n3653 ;
  assign n3656 = n3654 ^ n3650 ;
  assign n3661 = n3658 ^ n3656 ;
  assign n3649 = n3644 ^ n3643 ;
  assign n3662 = n3661 ^ n3649 ;
  assign n3741 = n3694 ^ n3662 ;
  assign n3764 = n3753 ^ n3741 ;
  assign n3765 = n3764 ^ n3607 ;
  assign n3280 = n3275 ^ n3273 ;
  assign n3281 = n3276 ^ n3274 ;
  assign n3282 = n3280 & n3281 ;
  assign n3284 = n3282 ^ n3278 ;
  assign n3289 = n3286 ^ n3284 ;
  assign n3277 = n3272 ^ n3271 ;
  assign n3290 = n3289 ^ n3277 ;
  assign n3248 = n3243 ^ n3241 ;
  assign n3249 = n3244 ^ n3242 ;
  assign n3250 = n3248 & n3249 ;
  assign n3252 = n3250 ^ n3246 ;
  assign n3257 = n3254 ^ n3252 ;
  assign n3245 = n3240 ^ n3239 ;
  assign n3258 = n3257 ^ n3245 ;
  assign n3337 = n3290 ^ n3258 ;
  assign n3360 = n3349 ^ n3337 ;
  assign n3361 = n3360 ^ n3203 ;
  assign n4236 = n3765 ^ n3361 ;
  assign n4327 = n4284 ^ n4236 ;
  assign n4328 = n4327 ^ n2862 ;
  assign n12827 = n8440 ^ n4328 ;
  assign n7813 = n7734 ^ n7726 ;
  assign n7814 = n7735 ^ n7727 ;
  assign n7826 = n7813 & n7814 ;
  assign n7811 = n7732 ^ n7724 ;
  assign n7812 = n7733 ^ n7725 ;
  assign n7825 = n7811 & n7812 ;
  assign n7830 = n7826 ^ n7825 ;
  assign n7809 = n7730 ^ n7722 ;
  assign n7810 = n7731 ^ n7723 ;
  assign n7819 = n7809 & n7810 ;
  assign n7807 = n7728 ^ n7720 ;
  assign n7808 = n7729 ^ n7721 ;
  assign n7818 = n7807 & n7808 ;
  assign n7823 = n7819 ^ n7818 ;
  assign n7844 = n7830 ^ n7823 ;
  assign n7854 = n7850 ^ n7844 ;
  assign n7855 = n7854 ^ n7804 ;
  assign n7878 = n7866 ^ n7855 ;
  assign n7739 = n7717 ^ n7708 ;
  assign n7879 = n7878 ^ n7739 ;
  assign n7409 = n7330 ^ n7322 ;
  assign n7410 = n7331 ^ n7323 ;
  assign n7422 = n7409 & n7410 ;
  assign n7407 = n7328 ^ n7320 ;
  assign n7408 = n7329 ^ n7321 ;
  assign n7421 = n7407 & n7408 ;
  assign n7426 = n7422 ^ n7421 ;
  assign n7405 = n7326 ^ n7318 ;
  assign n7406 = n7327 ^ n7319 ;
  assign n7415 = n7405 & n7406 ;
  assign n7403 = n7324 ^ n7316 ;
  assign n7404 = n7325 ^ n7317 ;
  assign n7414 = n7403 & n7404 ;
  assign n7419 = n7415 ^ n7414 ;
  assign n7440 = n7426 ^ n7419 ;
  assign n7450 = n7446 ^ n7440 ;
  assign n7451 = n7450 ^ n7400 ;
  assign n7474 = n7462 ^ n7451 ;
  assign n7335 = n7313 ^ n7304 ;
  assign n7475 = n7474 ^ n7335 ;
  assign n8349 = n7879 ^ n7475 ;
  assign n8441 = n8397 ^ n8349 ;
  assign n8442 = n8441 ^ n6976 ;
  assign n3701 = n3622 ^ n3614 ;
  assign n3702 = n3623 ^ n3615 ;
  assign n3714 = n3701 & n3702 ;
  assign n3699 = n3620 ^ n3612 ;
  assign n3700 = n3621 ^ n3613 ;
  assign n3713 = n3699 & n3700 ;
  assign n3718 = n3714 ^ n3713 ;
  assign n3697 = n3618 ^ n3610 ;
  assign n3698 = n3619 ^ n3611 ;
  assign n3707 = n3697 & n3698 ;
  assign n3695 = n3616 ^ n3608 ;
  assign n3696 = n3617 ^ n3609 ;
  assign n3706 = n3695 & n3696 ;
  assign n3711 = n3707 ^ n3706 ;
  assign n3732 = n3718 ^ n3711 ;
  assign n3742 = n3738 ^ n3732 ;
  assign n3743 = n3742 ^ n3692 ;
  assign n3766 = n3754 ^ n3743 ;
  assign n3627 = n3605 ^ n3596 ;
  assign n3767 = n3766 ^ n3627 ;
  assign n3297 = n3218 ^ n3210 ;
  assign n3298 = n3219 ^ n3211 ;
  assign n3310 = n3297 & n3298 ;
  assign n3295 = n3216 ^ n3208 ;
  assign n3296 = n3217 ^ n3209 ;
  assign n3309 = n3295 & n3296 ;
  assign n3314 = n3310 ^ n3309 ;
  assign n3293 = n3214 ^ n3206 ;
  assign n3294 = n3215 ^ n3207 ;
  assign n3303 = n3293 & n3294 ;
  assign n3291 = n3212 ^ n3204 ;
  assign n3292 = n3213 ^ n3205 ;
  assign n3302 = n3291 & n3292 ;
  assign n3307 = n3303 ^ n3302 ;
  assign n3328 = n3314 ^ n3307 ;
  assign n3338 = n3334 ^ n3328 ;
  assign n3339 = n3338 ^ n3288 ;
  assign n3362 = n3350 ^ n3339 ;
  assign n3223 = n3201 ^ n3192 ;
  assign n3363 = n3362 ^ n3223 ;
  assign n4237 = n3767 ^ n3363 ;
  assign n4329 = n4285 ^ n4237 ;
  assign n4330 = n4329 ^ n2864 ;
  assign n12828 = n8442 ^ n4330 ;
  assign n7827 = n7813 ^ n7811 ;
  assign n7828 = n7814 ^ n7812 ;
  assign n7829 = n7827 & n7828 ;
  assign n7831 = n7829 ^ n7825 ;
  assign n7820 = n7809 ^ n7807 ;
  assign n7821 = n7810 ^ n7808 ;
  assign n7822 = n7820 & n7821 ;
  assign n7824 = n7822 ^ n7818 ;
  assign n7845 = n7831 ^ n7824 ;
  assign n7856 = n7851 ^ n7845 ;
  assign n7857 = n7856 ^ n7806 ;
  assign n7880 = n7867 ^ n7857 ;
  assign n7740 = n7719 ^ n7709 ;
  assign n7881 = n7880 ^ n7740 ;
  assign n7423 = n7409 ^ n7407 ;
  assign n7424 = n7410 ^ n7408 ;
  assign n7425 = n7423 & n7424 ;
  assign n7427 = n7425 ^ n7421 ;
  assign n7416 = n7405 ^ n7403 ;
  assign n7417 = n7406 ^ n7404 ;
  assign n7418 = n7416 & n7417 ;
  assign n7420 = n7418 ^ n7414 ;
  assign n7441 = n7427 ^ n7420 ;
  assign n7452 = n7447 ^ n7441 ;
  assign n7453 = n7452 ^ n7402 ;
  assign n7476 = n7463 ^ n7453 ;
  assign n7336 = n7315 ^ n7305 ;
  assign n7477 = n7476 ^ n7336 ;
  assign n8350 = n7881 ^ n7477 ;
  assign n8443 = n8398 ^ n8350 ;
  assign n8444 = n8443 ^ n6978 ;
  assign n3715 = n3701 ^ n3699 ;
  assign n3716 = n3702 ^ n3700 ;
  assign n3717 = n3715 & n3716 ;
  assign n3719 = n3717 ^ n3713 ;
  assign n3708 = n3697 ^ n3695 ;
  assign n3709 = n3698 ^ n3696 ;
  assign n3710 = n3708 & n3709 ;
  assign n3712 = n3710 ^ n3706 ;
  assign n3733 = n3719 ^ n3712 ;
  assign n3744 = n3739 ^ n3733 ;
  assign n3745 = n3744 ^ n3694 ;
  assign n3768 = n3755 ^ n3745 ;
  assign n3628 = n3607 ^ n3597 ;
  assign n3769 = n3768 ^ n3628 ;
  assign n3311 = n3297 ^ n3295 ;
  assign n3312 = n3298 ^ n3296 ;
  assign n3313 = n3311 & n3312 ;
  assign n3315 = n3313 ^ n3309 ;
  assign n3304 = n3293 ^ n3291 ;
  assign n3305 = n3294 ^ n3292 ;
  assign n3306 = n3304 & n3305 ;
  assign n3308 = n3306 ^ n3302 ;
  assign n3329 = n3315 ^ n3308 ;
  assign n3340 = n3335 ^ n3329 ;
  assign n3341 = n3340 ^ n3290 ;
  assign n3364 = n3351 ^ n3341 ;
  assign n3224 = n3203 ^ n3193 ;
  assign n3365 = n3364 ^ n3224 ;
  assign n4238 = n3769 ^ n3365 ;
  assign n4331 = n4286 ^ n4238 ;
  assign n4332 = n4331 ^ n2866 ;
  assign n12829 = n8444 ^ n4332 ;
  assign n7834 = n7813 ^ n7809 ;
  assign n7835 = n7814 ^ n7810 ;
  assign n7838 = n7834 & n7835 ;
  assign n7832 = n7811 ^ n7807 ;
  assign n7833 = n7812 ^ n7808 ;
  assign n7837 = n7832 & n7833 ;
  assign n7842 = n7838 ^ n7837 ;
  assign n7846 = n7844 ^ n7842 ;
  assign n7847 = n7846 ^ n7831 ;
  assign n7858 = n7852 ^ n7847 ;
  assign n7816 = n7806 ^ n7801 ;
  assign n7859 = n7858 ^ n7816 ;
  assign n7882 = n7868 ^ n7859 ;
  assign n7737 = n7719 ^ n7713 ;
  assign n7741 = n7737 ^ n7710 ;
  assign n7883 = n7882 ^ n7741 ;
  assign n7430 = n7409 ^ n7405 ;
  assign n7431 = n7410 ^ n7406 ;
  assign n7434 = n7430 & n7431 ;
  assign n7428 = n7407 ^ n7403 ;
  assign n7429 = n7408 ^ n7404 ;
  assign n7433 = n7428 & n7429 ;
  assign n7438 = n7434 ^ n7433 ;
  assign n7442 = n7440 ^ n7438 ;
  assign n7443 = n7442 ^ n7427 ;
  assign n7454 = n7448 ^ n7443 ;
  assign n7412 = n7402 ^ n7397 ;
  assign n7455 = n7454 ^ n7412 ;
  assign n7478 = n7464 ^ n7455 ;
  assign n7333 = n7315 ^ n7309 ;
  assign n7337 = n7333 ^ n7306 ;
  assign n7479 = n7478 ^ n7337 ;
  assign n8351 = n7883 ^ n7479 ;
  assign n8445 = n8399 ^ n8351 ;
  assign n8446 = n8445 ^ n6980 ;
  assign n3722 = n3701 ^ n3697 ;
  assign n3723 = n3702 ^ n3698 ;
  assign n3726 = n3722 & n3723 ;
  assign n3720 = n3699 ^ n3695 ;
  assign n3721 = n3700 ^ n3696 ;
  assign n3725 = n3720 & n3721 ;
  assign n3730 = n3726 ^ n3725 ;
  assign n3734 = n3732 ^ n3730 ;
  assign n3735 = n3734 ^ n3719 ;
  assign n3746 = n3740 ^ n3735 ;
  assign n3704 = n3694 ^ n3689 ;
  assign n3747 = n3746 ^ n3704 ;
  assign n3770 = n3756 ^ n3747 ;
  assign n3625 = n3607 ^ n3601 ;
  assign n3629 = n3625 ^ n3598 ;
  assign n3771 = n3770 ^ n3629 ;
  assign n3318 = n3297 ^ n3293 ;
  assign n3319 = n3298 ^ n3294 ;
  assign n3322 = n3318 & n3319 ;
  assign n3316 = n3295 ^ n3291 ;
  assign n3317 = n3296 ^ n3292 ;
  assign n3321 = n3316 & n3317 ;
  assign n3326 = n3322 ^ n3321 ;
  assign n3330 = n3328 ^ n3326 ;
  assign n3331 = n3330 ^ n3315 ;
  assign n3342 = n3336 ^ n3331 ;
  assign n3300 = n3290 ^ n3285 ;
  assign n3343 = n3342 ^ n3300 ;
  assign n3366 = n3352 ^ n3343 ;
  assign n3221 = n3203 ^ n3197 ;
  assign n3225 = n3221 ^ n3194 ;
  assign n3367 = n3366 ^ n3225 ;
  assign n4239 = n3771 ^ n3367 ;
  assign n4333 = n4287 ^ n4239 ;
  assign n4334 = n4333 ^ n2868 ;
  assign n12830 = n8446 ^ n4334 ;
  assign n7839 = n7834 ^ n7832 ;
  assign n7840 = n7835 ^ n7833 ;
  assign n7841 = n7839 & n7840 ;
  assign n7843 = n7841 ^ n7837 ;
  assign n7848 = n7845 ^ n7843 ;
  assign n7836 = n7831 ^ n7830 ;
  assign n7849 = n7848 ^ n7836 ;
  assign n7860 = n7853 ^ n7849 ;
  assign n7815 = n7806 ^ n7804 ;
  assign n7817 = n7815 ^ n7802 ;
  assign n7861 = n7860 ^ n7817 ;
  assign n7884 = n7869 ^ n7861 ;
  assign n7736 = n7719 ^ n7717 ;
  assign n7738 = n7736 ^ n7715 ;
  assign n7742 = n7738 ^ n7711 ;
  assign n7885 = n7884 ^ n7742 ;
  assign n7435 = n7430 ^ n7428 ;
  assign n7436 = n7431 ^ n7429 ;
  assign n7437 = n7435 & n7436 ;
  assign n7439 = n7437 ^ n7433 ;
  assign n7444 = n7441 ^ n7439 ;
  assign n7432 = n7427 ^ n7426 ;
  assign n7445 = n7444 ^ n7432 ;
  assign n7456 = n7449 ^ n7445 ;
  assign n7411 = n7402 ^ n7400 ;
  assign n7413 = n7411 ^ n7398 ;
  assign n7457 = n7456 ^ n7413 ;
  assign n7480 = n7465 ^ n7457 ;
  assign n7332 = n7315 ^ n7313 ;
  assign n7334 = n7332 ^ n7311 ;
  assign n7338 = n7334 ^ n7307 ;
  assign n7481 = n7480 ^ n7338 ;
  assign n8352 = n7885 ^ n7481 ;
  assign n8447 = n8400 ^ n8352 ;
  assign n8448 = n8447 ^ n6982 ;
  assign n3727 = n3722 ^ n3720 ;
  assign n3728 = n3723 ^ n3721 ;
  assign n3729 = n3727 & n3728 ;
  assign n3731 = n3729 ^ n3725 ;
  assign n3736 = n3733 ^ n3731 ;
  assign n3724 = n3719 ^ n3718 ;
  assign n3737 = n3736 ^ n3724 ;
  assign n3748 = n3741 ^ n3737 ;
  assign n3703 = n3694 ^ n3692 ;
  assign n3705 = n3703 ^ n3690 ;
  assign n3749 = n3748 ^ n3705 ;
  assign n3772 = n3757 ^ n3749 ;
  assign n3624 = n3607 ^ n3605 ;
  assign n3626 = n3624 ^ n3603 ;
  assign n3630 = n3626 ^ n3599 ;
  assign n3773 = n3772 ^ n3630 ;
  assign n3323 = n3318 ^ n3316 ;
  assign n3324 = n3319 ^ n3317 ;
  assign n3325 = n3323 & n3324 ;
  assign n3327 = n3325 ^ n3321 ;
  assign n3332 = n3329 ^ n3327 ;
  assign n3320 = n3315 ^ n3314 ;
  assign n3333 = n3332 ^ n3320 ;
  assign n3344 = n3337 ^ n3333 ;
  assign n3299 = n3290 ^ n3288 ;
  assign n3301 = n3299 ^ n3286 ;
  assign n3345 = n3344 ^ n3301 ;
  assign n3368 = n3353 ^ n3345 ;
  assign n3220 = n3203 ^ n3201 ;
  assign n3222 = n3220 ^ n3199 ;
  assign n3226 = n3222 ^ n3195 ;
  assign n3369 = n3368 ^ n3226 ;
  assign n4240 = n3773 ^ n3369 ;
  assign n4335 = n4288 ^ n4240 ;
  assign n4336 = n4335 ^ n2870 ;
  assign n12831 = n8448 ^ n4336 ;
  assign n7916 = n7045 ^ n7013 ;
  assign n7917 = n7046 ^ n7014 ;
  assign n8092 = n7916 & n7917 ;
  assign n7914 = n7043 ^ n7011 ;
  assign n7915 = n7044 ^ n7012 ;
  assign n8091 = n7914 & n7915 ;
  assign n8096 = n8092 ^ n8091 ;
  assign n7912 = n7041 ^ n7009 ;
  assign n7913 = n7042 ^ n7010 ;
  assign n8085 = n7912 & n7913 ;
  assign n7910 = n7039 ^ n7007 ;
  assign n7911 = n7040 ^ n7008 ;
  assign n8084 = n7910 & n7911 ;
  assign n8089 = n8085 ^ n8084 ;
  assign n8110 = n8096 ^ n8089 ;
  assign n7908 = n7037 ^ n7005 ;
  assign n7909 = n7038 ^ n7006 ;
  assign n8060 = n7908 & n7909 ;
  assign n7906 = n7035 ^ n7003 ;
  assign n7907 = n7036 ^ n7004 ;
  assign n8059 = n7906 & n7907 ;
  assign n8064 = n8060 ^ n8059 ;
  assign n7904 = n7033 ^ n7001 ;
  assign n7905 = n7034 ^ n7002 ;
  assign n8053 = n7904 & n7905 ;
  assign n7902 = n7031 ^ n6999 ;
  assign n7903 = n7032 ^ n7000 ;
  assign n8052 = n7902 & n7903 ;
  assign n8057 = n8053 ^ n8052 ;
  assign n8078 = n8064 ^ n8057 ;
  assign n8159 = n8110 ^ n8078 ;
  assign n7900 = n7029 ^ n6997 ;
  assign n7901 = n7030 ^ n6998 ;
  assign n7973 = n7900 & n7901 ;
  assign n7898 = n7027 ^ n6995 ;
  assign n7899 = n7028 ^ n6996 ;
  assign n7972 = n7898 & n7899 ;
  assign n7977 = n7973 ^ n7972 ;
  assign n7896 = n7025 ^ n6993 ;
  assign n7897 = n7026 ^ n6994 ;
  assign n7966 = n7896 & n7897 ;
  assign n7894 = n7023 ^ n6991 ;
  assign n7895 = n7024 ^ n6992 ;
  assign n7965 = n7894 & n7895 ;
  assign n7970 = n7966 ^ n7965 ;
  assign n7991 = n7977 ^ n7970 ;
  assign n7892 = n7021 ^ n6989 ;
  assign n7893 = n7022 ^ n6990 ;
  assign n7941 = n7892 & n7893 ;
  assign n7890 = n7019 ^ n6987 ;
  assign n7891 = n7020 ^ n6988 ;
  assign n7940 = n7890 & n7891 ;
  assign n7945 = n7941 ^ n7940 ;
  assign n7888 = n7017 ^ n6985 ;
  assign n7889 = n7018 ^ n6986 ;
  assign n7934 = n7888 & n7889 ;
  assign n7886 = n7015 ^ n6983 ;
  assign n7887 = n7016 ^ n6984 ;
  assign n7933 = n7886 & n7887 ;
  assign n7938 = n7934 ^ n7933 ;
  assign n7959 = n7945 ^ n7938 ;
  assign n8040 = n7991 ^ n7959 ;
  assign n8313 = n8159 ^ n8040 ;
  assign n8353 = n8337 ^ n8313 ;
  assign n8354 = n8353 ^ n7871 ;
  assign n8449 = n8401 ^ n8354 ;
  assign n7062 = n6968 ^ n6935 ;
  assign n8450 = n8449 ^ n7062 ;
  assign n3804 = n2933 ^ n2901 ;
  assign n3805 = n2934 ^ n2902 ;
  assign n3980 = n3804 & n3805 ;
  assign n3802 = n2931 ^ n2899 ;
  assign n3803 = n2932 ^ n2900 ;
  assign n3979 = n3802 & n3803 ;
  assign n3984 = n3980 ^ n3979 ;
  assign n3800 = n2929 ^ n2897 ;
  assign n3801 = n2930 ^ n2898 ;
  assign n3973 = n3800 & n3801 ;
  assign n3798 = n2927 ^ n2895 ;
  assign n3799 = n2928 ^ n2896 ;
  assign n3972 = n3798 & n3799 ;
  assign n3977 = n3973 ^ n3972 ;
  assign n3998 = n3984 ^ n3977 ;
  assign n3796 = n2925 ^ n2893 ;
  assign n3797 = n2926 ^ n2894 ;
  assign n3948 = n3796 & n3797 ;
  assign n3794 = n2923 ^ n2891 ;
  assign n3795 = n2924 ^ n2892 ;
  assign n3947 = n3794 & n3795 ;
  assign n3952 = n3948 ^ n3947 ;
  assign n3792 = n2921 ^ n2889 ;
  assign n3793 = n2922 ^ n2890 ;
  assign n3941 = n3792 & n3793 ;
  assign n3790 = n2919 ^ n2887 ;
  assign n3791 = n2920 ^ n2888 ;
  assign n3940 = n3790 & n3791 ;
  assign n3945 = n3941 ^ n3940 ;
  assign n3966 = n3952 ^ n3945 ;
  assign n4047 = n3998 ^ n3966 ;
  assign n3788 = n2917 ^ n2885 ;
  assign n3789 = n2918 ^ n2886 ;
  assign n3861 = n3788 & n3789 ;
  assign n3786 = n2915 ^ n2883 ;
  assign n3787 = n2916 ^ n2884 ;
  assign n3860 = n3786 & n3787 ;
  assign n3865 = n3861 ^ n3860 ;
  assign n3784 = n2913 ^ n2881 ;
  assign n3785 = n2914 ^ n2882 ;
  assign n3854 = n3784 & n3785 ;
  assign n3782 = n2911 ^ n2879 ;
  assign n3783 = n2912 ^ n2880 ;
  assign n3853 = n3782 & n3783 ;
  assign n3858 = n3854 ^ n3853 ;
  assign n3879 = n3865 ^ n3858 ;
  assign n3780 = n2909 ^ n2877 ;
  assign n3781 = n2910 ^ n2878 ;
  assign n3829 = n3780 & n3781 ;
  assign n3778 = n2907 ^ n2875 ;
  assign n3779 = n2908 ^ n2876 ;
  assign n3828 = n3778 & n3779 ;
  assign n3833 = n3829 ^ n3828 ;
  assign n3776 = n2905 ^ n2873 ;
  assign n3777 = n2906 ^ n2874 ;
  assign n3822 = n3776 & n3777 ;
  assign n3774 = n2903 ^ n2871 ;
  assign n3775 = n2904 ^ n2872 ;
  assign n3821 = n3774 & n3775 ;
  assign n3826 = n3822 ^ n3821 ;
  assign n3847 = n3833 ^ n3826 ;
  assign n3928 = n3879 ^ n3847 ;
  assign n4201 = n4047 ^ n3928 ;
  assign n4241 = n4225 ^ n4201 ;
  assign n4242 = n4241 ^ n3759 ;
  assign n4337 = n4289 ^ n4242 ;
  assign n2950 = n2856 ^ n2823 ;
  assign n4338 = n4337 ^ n2950 ;
  assign n12832 = n8450 ^ n4338 ;
  assign n8093 = n7916 ^ n7914 ;
  assign n8094 = n7917 ^ n7915 ;
  assign n8095 = n8093 & n8094 ;
  assign n8097 = n8095 ^ n8091 ;
  assign n8086 = n7912 ^ n7910 ;
  assign n8087 = n7913 ^ n7911 ;
  assign n8088 = n8086 & n8087 ;
  assign n8090 = n8088 ^ n8084 ;
  assign n8111 = n8097 ^ n8090 ;
  assign n8061 = n7908 ^ n7906 ;
  assign n8062 = n7909 ^ n7907 ;
  assign n8063 = n8061 & n8062 ;
  assign n8065 = n8063 ^ n8059 ;
  assign n8054 = n7904 ^ n7902 ;
  assign n8055 = n7905 ^ n7903 ;
  assign n8056 = n8054 & n8055 ;
  assign n8058 = n8056 ^ n8052 ;
  assign n8079 = n8065 ^ n8058 ;
  assign n8160 = n8111 ^ n8079 ;
  assign n7974 = n7900 ^ n7898 ;
  assign n7975 = n7901 ^ n7899 ;
  assign n7976 = n7974 & n7975 ;
  assign n7978 = n7976 ^ n7972 ;
  assign n7967 = n7896 ^ n7894 ;
  assign n7968 = n7897 ^ n7895 ;
  assign n7969 = n7967 & n7968 ;
  assign n7971 = n7969 ^ n7965 ;
  assign n7992 = n7978 ^ n7971 ;
  assign n7942 = n7892 ^ n7890 ;
  assign n7943 = n7893 ^ n7891 ;
  assign n7944 = n7942 & n7943 ;
  assign n7946 = n7944 ^ n7940 ;
  assign n7935 = n7888 ^ n7886 ;
  assign n7936 = n7889 ^ n7887 ;
  assign n7937 = n7935 & n7936 ;
  assign n7939 = n7937 ^ n7933 ;
  assign n7960 = n7946 ^ n7939 ;
  assign n8041 = n7992 ^ n7960 ;
  assign n8314 = n8160 ^ n8041 ;
  assign n8355 = n8338 ^ n8314 ;
  assign n8356 = n8355 ^ n7873 ;
  assign n8451 = n8402 ^ n8356 ;
  assign n7063 = n6970 ^ n6936 ;
  assign n8452 = n8451 ^ n7063 ;
  assign n3981 = n3804 ^ n3802 ;
  assign n3982 = n3805 ^ n3803 ;
  assign n3983 = n3981 & n3982 ;
  assign n3985 = n3983 ^ n3979 ;
  assign n3974 = n3800 ^ n3798 ;
  assign n3975 = n3801 ^ n3799 ;
  assign n3976 = n3974 & n3975 ;
  assign n3978 = n3976 ^ n3972 ;
  assign n3999 = n3985 ^ n3978 ;
  assign n3949 = n3796 ^ n3794 ;
  assign n3950 = n3797 ^ n3795 ;
  assign n3951 = n3949 & n3950 ;
  assign n3953 = n3951 ^ n3947 ;
  assign n3942 = n3792 ^ n3790 ;
  assign n3943 = n3793 ^ n3791 ;
  assign n3944 = n3942 & n3943 ;
  assign n3946 = n3944 ^ n3940 ;
  assign n3967 = n3953 ^ n3946 ;
  assign n4048 = n3999 ^ n3967 ;
  assign n3862 = n3788 ^ n3786 ;
  assign n3863 = n3789 ^ n3787 ;
  assign n3864 = n3862 & n3863 ;
  assign n3866 = n3864 ^ n3860 ;
  assign n3855 = n3784 ^ n3782 ;
  assign n3856 = n3785 ^ n3783 ;
  assign n3857 = n3855 & n3856 ;
  assign n3859 = n3857 ^ n3853 ;
  assign n3880 = n3866 ^ n3859 ;
  assign n3830 = n3780 ^ n3778 ;
  assign n3831 = n3781 ^ n3779 ;
  assign n3832 = n3830 & n3831 ;
  assign n3834 = n3832 ^ n3828 ;
  assign n3823 = n3776 ^ n3774 ;
  assign n3824 = n3777 ^ n3775 ;
  assign n3825 = n3823 & n3824 ;
  assign n3827 = n3825 ^ n3821 ;
  assign n3848 = n3834 ^ n3827 ;
  assign n3929 = n3880 ^ n3848 ;
  assign n4202 = n4048 ^ n3929 ;
  assign n4243 = n4226 ^ n4202 ;
  assign n4244 = n4243 ^ n3761 ;
  assign n4339 = n4290 ^ n4244 ;
  assign n2951 = n2858 ^ n2824 ;
  assign n4340 = n4339 ^ n2951 ;
  assign n12833 = n8452 ^ n4340 ;
  assign n8100 = n7916 ^ n7912 ;
  assign n8101 = n7917 ^ n7913 ;
  assign n8104 = n8100 & n8101 ;
  assign n8098 = n7914 ^ n7910 ;
  assign n8099 = n7915 ^ n7911 ;
  assign n8103 = n8098 & n8099 ;
  assign n8108 = n8104 ^ n8103 ;
  assign n8112 = n8110 ^ n8108 ;
  assign n8113 = n8112 ^ n8097 ;
  assign n8068 = n7908 ^ n7904 ;
  assign n8069 = n7909 ^ n7905 ;
  assign n8072 = n8068 & n8069 ;
  assign n8066 = n7906 ^ n7902 ;
  assign n8067 = n7907 ^ n7903 ;
  assign n8071 = n8066 & n8067 ;
  assign n8076 = n8072 ^ n8071 ;
  assign n8080 = n8078 ^ n8076 ;
  assign n8081 = n8080 ^ n8065 ;
  assign n8161 = n8113 ^ n8081 ;
  assign n7981 = n7900 ^ n7896 ;
  assign n7982 = n7901 ^ n7897 ;
  assign n7985 = n7981 & n7982 ;
  assign n7979 = n7898 ^ n7894 ;
  assign n7980 = n7899 ^ n7895 ;
  assign n7984 = n7979 & n7980 ;
  assign n7989 = n7985 ^ n7984 ;
  assign n7993 = n7991 ^ n7989 ;
  assign n7994 = n7993 ^ n7978 ;
  assign n7949 = n7892 ^ n7888 ;
  assign n7950 = n7893 ^ n7889 ;
  assign n7953 = n7949 & n7950 ;
  assign n7947 = n7890 ^ n7886 ;
  assign n7948 = n7891 ^ n7887 ;
  assign n7952 = n7947 & n7948 ;
  assign n7957 = n7953 ^ n7952 ;
  assign n7961 = n7959 ^ n7957 ;
  assign n7962 = n7961 ^ n7946 ;
  assign n8042 = n7994 ^ n7962 ;
  assign n8315 = n8161 ^ n8042 ;
  assign n8357 = n8339 ^ n8315 ;
  assign n8358 = n8357 ^ n7875 ;
  assign n8453 = n8403 ^ n8358 ;
  assign n7064 = n6972 ^ n6937 ;
  assign n8454 = n8453 ^ n7064 ;
  assign n3988 = n3804 ^ n3800 ;
  assign n3989 = n3805 ^ n3801 ;
  assign n3992 = n3988 & n3989 ;
  assign n3986 = n3802 ^ n3798 ;
  assign n3987 = n3803 ^ n3799 ;
  assign n3991 = n3986 & n3987 ;
  assign n3996 = n3992 ^ n3991 ;
  assign n4000 = n3998 ^ n3996 ;
  assign n4001 = n4000 ^ n3985 ;
  assign n3956 = n3796 ^ n3792 ;
  assign n3957 = n3797 ^ n3793 ;
  assign n3960 = n3956 & n3957 ;
  assign n3954 = n3794 ^ n3790 ;
  assign n3955 = n3795 ^ n3791 ;
  assign n3959 = n3954 & n3955 ;
  assign n3964 = n3960 ^ n3959 ;
  assign n3968 = n3966 ^ n3964 ;
  assign n3969 = n3968 ^ n3953 ;
  assign n4049 = n4001 ^ n3969 ;
  assign n3869 = n3788 ^ n3784 ;
  assign n3870 = n3789 ^ n3785 ;
  assign n3873 = n3869 & n3870 ;
  assign n3867 = n3786 ^ n3782 ;
  assign n3868 = n3787 ^ n3783 ;
  assign n3872 = n3867 & n3868 ;
  assign n3877 = n3873 ^ n3872 ;
  assign n3881 = n3879 ^ n3877 ;
  assign n3882 = n3881 ^ n3866 ;
  assign n3837 = n3780 ^ n3776 ;
  assign n3838 = n3781 ^ n3777 ;
  assign n3841 = n3837 & n3838 ;
  assign n3835 = n3778 ^ n3774 ;
  assign n3836 = n3779 ^ n3775 ;
  assign n3840 = n3835 & n3836 ;
  assign n3845 = n3841 ^ n3840 ;
  assign n3849 = n3847 ^ n3845 ;
  assign n3850 = n3849 ^ n3834 ;
  assign n3930 = n3882 ^ n3850 ;
  assign n4203 = n4049 ^ n3930 ;
  assign n4245 = n4227 ^ n4203 ;
  assign n4246 = n4245 ^ n3763 ;
  assign n4341 = n4291 ^ n4246 ;
  assign n2952 = n2860 ^ n2825 ;
  assign n4342 = n4341 ^ n2952 ;
  assign n12834 = n8454 ^ n4342 ;
  assign n8105 = n8100 ^ n8098 ;
  assign n8106 = n8101 ^ n8099 ;
  assign n8107 = n8105 & n8106 ;
  assign n8109 = n8107 ^ n8103 ;
  assign n8114 = n8111 ^ n8109 ;
  assign n8102 = n8097 ^ n8096 ;
  assign n8115 = n8114 ^ n8102 ;
  assign n8073 = n8068 ^ n8066 ;
  assign n8074 = n8069 ^ n8067 ;
  assign n8075 = n8073 & n8074 ;
  assign n8077 = n8075 ^ n8071 ;
  assign n8082 = n8079 ^ n8077 ;
  assign n8070 = n8065 ^ n8064 ;
  assign n8083 = n8082 ^ n8070 ;
  assign n8162 = n8115 ^ n8083 ;
  assign n7986 = n7981 ^ n7979 ;
  assign n7987 = n7982 ^ n7980 ;
  assign n7988 = n7986 & n7987 ;
  assign n7990 = n7988 ^ n7984 ;
  assign n7995 = n7992 ^ n7990 ;
  assign n7983 = n7978 ^ n7977 ;
  assign n7996 = n7995 ^ n7983 ;
  assign n7954 = n7949 ^ n7947 ;
  assign n7955 = n7950 ^ n7948 ;
  assign n7956 = n7954 & n7955 ;
  assign n7958 = n7956 ^ n7952 ;
  assign n7963 = n7960 ^ n7958 ;
  assign n7951 = n7946 ^ n7945 ;
  assign n7964 = n7963 ^ n7951 ;
  assign n8043 = n7996 ^ n7964 ;
  assign n8316 = n8162 ^ n8043 ;
  assign n8359 = n8340 ^ n8316 ;
  assign n8360 = n8359 ^ n7877 ;
  assign n8455 = n8404 ^ n8360 ;
  assign n7065 = n6974 ^ n6938 ;
  assign n8456 = n8455 ^ n7065 ;
  assign n3993 = n3988 ^ n3986 ;
  assign n3994 = n3989 ^ n3987 ;
  assign n3995 = n3993 & n3994 ;
  assign n3997 = n3995 ^ n3991 ;
  assign n4002 = n3999 ^ n3997 ;
  assign n3990 = n3985 ^ n3984 ;
  assign n4003 = n4002 ^ n3990 ;
  assign n3961 = n3956 ^ n3954 ;
  assign n3962 = n3957 ^ n3955 ;
  assign n3963 = n3961 & n3962 ;
  assign n3965 = n3963 ^ n3959 ;
  assign n3970 = n3967 ^ n3965 ;
  assign n3958 = n3953 ^ n3952 ;
  assign n3971 = n3970 ^ n3958 ;
  assign n4050 = n4003 ^ n3971 ;
  assign n3874 = n3869 ^ n3867 ;
  assign n3875 = n3870 ^ n3868 ;
  assign n3876 = n3874 & n3875 ;
  assign n3878 = n3876 ^ n3872 ;
  assign n3883 = n3880 ^ n3878 ;
  assign n3871 = n3866 ^ n3865 ;
  assign n3884 = n3883 ^ n3871 ;
  assign n3842 = n3837 ^ n3835 ;
  assign n3843 = n3838 ^ n3836 ;
  assign n3844 = n3842 & n3843 ;
  assign n3846 = n3844 ^ n3840 ;
  assign n3851 = n3848 ^ n3846 ;
  assign n3839 = n3834 ^ n3833 ;
  assign n3852 = n3851 ^ n3839 ;
  assign n3931 = n3884 ^ n3852 ;
  assign n4204 = n4050 ^ n3931 ;
  assign n4247 = n4228 ^ n4204 ;
  assign n4248 = n4247 ^ n3765 ;
  assign n4343 = n4292 ^ n4248 ;
  assign n2953 = n2862 ^ n2826 ;
  assign n4344 = n4343 ^ n2953 ;
  assign n12835 = n8456 ^ n4344 ;
  assign n8122 = n7916 ^ n7908 ;
  assign n8123 = n7917 ^ n7909 ;
  assign n8135 = n8122 & n8123 ;
  assign n8120 = n7914 ^ n7906 ;
  assign n8121 = n7915 ^ n7907 ;
  assign n8134 = n8120 & n8121 ;
  assign n8139 = n8135 ^ n8134 ;
  assign n8118 = n7912 ^ n7904 ;
  assign n8119 = n7913 ^ n7905 ;
  assign n8128 = n8118 & n8119 ;
  assign n8116 = n7910 ^ n7902 ;
  assign n8117 = n7911 ^ n7903 ;
  assign n8127 = n8116 & n8117 ;
  assign n8132 = n8128 ^ n8127 ;
  assign n8153 = n8139 ^ n8132 ;
  assign n8163 = n8159 ^ n8153 ;
  assign n8164 = n8163 ^ n8113 ;
  assign n8003 = n7900 ^ n7892 ;
  assign n8004 = n7901 ^ n7893 ;
  assign n8016 = n8003 & n8004 ;
  assign n8001 = n7898 ^ n7890 ;
  assign n8002 = n7899 ^ n7891 ;
  assign n8015 = n8001 & n8002 ;
  assign n8020 = n8016 ^ n8015 ;
  assign n7999 = n7896 ^ n7888 ;
  assign n8000 = n7897 ^ n7889 ;
  assign n8009 = n7999 & n8000 ;
  assign n7997 = n7894 ^ n7886 ;
  assign n7998 = n7895 ^ n7887 ;
  assign n8008 = n7997 & n7998 ;
  assign n8013 = n8009 ^ n8008 ;
  assign n8034 = n8020 ^ n8013 ;
  assign n8044 = n8040 ^ n8034 ;
  assign n8045 = n8044 ^ n7994 ;
  assign n8317 = n8164 ^ n8045 ;
  assign n8361 = n8341 ^ n8317 ;
  assign n8362 = n8361 ^ n7879 ;
  assign n8457 = n8405 ^ n8362 ;
  assign n7066 = n6976 ^ n6939 ;
  assign n8458 = n8457 ^ n7066 ;
  assign n4010 = n3804 ^ n3796 ;
  assign n4011 = n3805 ^ n3797 ;
  assign n4023 = n4010 & n4011 ;
  assign n4008 = n3802 ^ n3794 ;
  assign n4009 = n3803 ^ n3795 ;
  assign n4022 = n4008 & n4009 ;
  assign n4027 = n4023 ^ n4022 ;
  assign n4006 = n3800 ^ n3792 ;
  assign n4007 = n3801 ^ n3793 ;
  assign n4016 = n4006 & n4007 ;
  assign n4004 = n3798 ^ n3790 ;
  assign n4005 = n3799 ^ n3791 ;
  assign n4015 = n4004 & n4005 ;
  assign n4020 = n4016 ^ n4015 ;
  assign n4041 = n4027 ^ n4020 ;
  assign n4051 = n4047 ^ n4041 ;
  assign n4052 = n4051 ^ n4001 ;
  assign n3891 = n3788 ^ n3780 ;
  assign n3892 = n3789 ^ n3781 ;
  assign n3904 = n3891 & n3892 ;
  assign n3889 = n3786 ^ n3778 ;
  assign n3890 = n3787 ^ n3779 ;
  assign n3903 = n3889 & n3890 ;
  assign n3908 = n3904 ^ n3903 ;
  assign n3887 = n3784 ^ n3776 ;
  assign n3888 = n3785 ^ n3777 ;
  assign n3897 = n3887 & n3888 ;
  assign n3885 = n3782 ^ n3774 ;
  assign n3886 = n3783 ^ n3775 ;
  assign n3896 = n3885 & n3886 ;
  assign n3901 = n3897 ^ n3896 ;
  assign n3922 = n3908 ^ n3901 ;
  assign n3932 = n3928 ^ n3922 ;
  assign n3933 = n3932 ^ n3882 ;
  assign n4205 = n4052 ^ n3933 ;
  assign n4249 = n4229 ^ n4205 ;
  assign n4250 = n4249 ^ n3767 ;
  assign n4345 = n4293 ^ n4250 ;
  assign n2954 = n2864 ^ n2827 ;
  assign n4346 = n4345 ^ n2954 ;
  assign n12836 = n8458 ^ n4346 ;
  assign n8136 = n8122 ^ n8120 ;
  assign n8137 = n8123 ^ n8121 ;
  assign n8138 = n8136 & n8137 ;
  assign n8140 = n8138 ^ n8134 ;
  assign n8129 = n8118 ^ n8116 ;
  assign n8130 = n8119 ^ n8117 ;
  assign n8131 = n8129 & n8130 ;
  assign n8133 = n8131 ^ n8127 ;
  assign n8154 = n8140 ^ n8133 ;
  assign n8165 = n8160 ^ n8154 ;
  assign n8166 = n8165 ^ n8115 ;
  assign n8017 = n8003 ^ n8001 ;
  assign n8018 = n8004 ^ n8002 ;
  assign n8019 = n8017 & n8018 ;
  assign n8021 = n8019 ^ n8015 ;
  assign n8010 = n7999 ^ n7997 ;
  assign n8011 = n8000 ^ n7998 ;
  assign n8012 = n8010 & n8011 ;
  assign n8014 = n8012 ^ n8008 ;
  assign n8035 = n8021 ^ n8014 ;
  assign n8046 = n8041 ^ n8035 ;
  assign n8047 = n8046 ^ n7996 ;
  assign n8318 = n8166 ^ n8047 ;
  assign n8363 = n8342 ^ n8318 ;
  assign n8364 = n8363 ^ n7881 ;
  assign n8459 = n8406 ^ n8364 ;
  assign n7067 = n6978 ^ n6940 ;
  assign n8460 = n8459 ^ n7067 ;
  assign n4024 = n4010 ^ n4008 ;
  assign n4025 = n4011 ^ n4009 ;
  assign n4026 = n4024 & n4025 ;
  assign n4028 = n4026 ^ n4022 ;
  assign n4017 = n4006 ^ n4004 ;
  assign n4018 = n4007 ^ n4005 ;
  assign n4019 = n4017 & n4018 ;
  assign n4021 = n4019 ^ n4015 ;
  assign n4042 = n4028 ^ n4021 ;
  assign n4053 = n4048 ^ n4042 ;
  assign n4054 = n4053 ^ n4003 ;
  assign n3905 = n3891 ^ n3889 ;
  assign n3906 = n3892 ^ n3890 ;
  assign n3907 = n3905 & n3906 ;
  assign n3909 = n3907 ^ n3903 ;
  assign n3898 = n3887 ^ n3885 ;
  assign n3899 = n3888 ^ n3886 ;
  assign n3900 = n3898 & n3899 ;
  assign n3902 = n3900 ^ n3896 ;
  assign n3923 = n3909 ^ n3902 ;
  assign n3934 = n3929 ^ n3923 ;
  assign n3935 = n3934 ^ n3884 ;
  assign n4206 = n4054 ^ n3935 ;
  assign n4251 = n4230 ^ n4206 ;
  assign n4252 = n4251 ^ n3769 ;
  assign n4347 = n4294 ^ n4252 ;
  assign n2955 = n2866 ^ n2828 ;
  assign n4348 = n4347 ^ n2955 ;
  assign n12837 = n8460 ^ n4348 ;
  assign n8143 = n8122 ^ n8118 ;
  assign n8144 = n8123 ^ n8119 ;
  assign n8147 = n8143 & n8144 ;
  assign n8141 = n8120 ^ n8116 ;
  assign n8142 = n8121 ^ n8117 ;
  assign n8146 = n8141 & n8142 ;
  assign n8151 = n8147 ^ n8146 ;
  assign n8155 = n8153 ^ n8151 ;
  assign n8156 = n8155 ^ n8140 ;
  assign n8167 = n8161 ^ n8156 ;
  assign n8125 = n8115 ^ n8110 ;
  assign n8168 = n8167 ^ n8125 ;
  assign n8024 = n8003 ^ n7999 ;
  assign n8025 = n8004 ^ n8000 ;
  assign n8028 = n8024 & n8025 ;
  assign n8022 = n8001 ^ n7997 ;
  assign n8023 = n8002 ^ n7998 ;
  assign n8027 = n8022 & n8023 ;
  assign n8032 = n8028 ^ n8027 ;
  assign n8036 = n8034 ^ n8032 ;
  assign n8037 = n8036 ^ n8021 ;
  assign n8048 = n8042 ^ n8037 ;
  assign n8006 = n7996 ^ n7991 ;
  assign n8049 = n8048 ^ n8006 ;
  assign n8319 = n8168 ^ n8049 ;
  assign n8365 = n8343 ^ n8319 ;
  assign n8366 = n8365 ^ n7883 ;
  assign n8461 = n8407 ^ n8366 ;
  assign n7068 = n6980 ^ n6941 ;
  assign n8462 = n8461 ^ n7068 ;
  assign n4031 = n4010 ^ n4006 ;
  assign n4032 = n4011 ^ n4007 ;
  assign n4035 = n4031 & n4032 ;
  assign n4029 = n4008 ^ n4004 ;
  assign n4030 = n4009 ^ n4005 ;
  assign n4034 = n4029 & n4030 ;
  assign n4039 = n4035 ^ n4034 ;
  assign n4043 = n4041 ^ n4039 ;
  assign n4044 = n4043 ^ n4028 ;
  assign n4055 = n4049 ^ n4044 ;
  assign n4013 = n4003 ^ n3998 ;
  assign n4056 = n4055 ^ n4013 ;
  assign n3912 = n3891 ^ n3887 ;
  assign n3913 = n3892 ^ n3888 ;
  assign n3916 = n3912 & n3913 ;
  assign n3910 = n3889 ^ n3885 ;
  assign n3911 = n3890 ^ n3886 ;
  assign n3915 = n3910 & n3911 ;
  assign n3920 = n3916 ^ n3915 ;
  assign n3924 = n3922 ^ n3920 ;
  assign n3925 = n3924 ^ n3909 ;
  assign n3936 = n3930 ^ n3925 ;
  assign n3894 = n3884 ^ n3879 ;
  assign n3937 = n3936 ^ n3894 ;
  assign n4207 = n4056 ^ n3937 ;
  assign n4253 = n4231 ^ n4207 ;
  assign n4254 = n4253 ^ n3771 ;
  assign n4349 = n4295 ^ n4254 ;
  assign n2956 = n2868 ^ n2829 ;
  assign n4350 = n4349 ^ n2956 ;
  assign n12838 = n8462 ^ n4350 ;
  assign n8148 = n8143 ^ n8141 ;
  assign n8149 = n8144 ^ n8142 ;
  assign n8150 = n8148 & n8149 ;
  assign n8152 = n8150 ^ n8146 ;
  assign n8157 = n8154 ^ n8152 ;
  assign n8145 = n8140 ^ n8139 ;
  assign n8158 = n8157 ^ n8145 ;
  assign n8169 = n8162 ^ n8158 ;
  assign n8124 = n8115 ^ n8113 ;
  assign n8126 = n8124 ^ n8111 ;
  assign n8170 = n8169 ^ n8126 ;
  assign n8029 = n8024 ^ n8022 ;
  assign n8030 = n8025 ^ n8023 ;
  assign n8031 = n8029 & n8030 ;
  assign n8033 = n8031 ^ n8027 ;
  assign n8038 = n8035 ^ n8033 ;
  assign n8026 = n8021 ^ n8020 ;
  assign n8039 = n8038 ^ n8026 ;
  assign n8050 = n8043 ^ n8039 ;
  assign n8005 = n7996 ^ n7994 ;
  assign n8007 = n8005 ^ n7992 ;
  assign n8051 = n8050 ^ n8007 ;
  assign n8320 = n8170 ^ n8051 ;
  assign n8367 = n8344 ^ n8320 ;
  assign n8368 = n8367 ^ n7885 ;
  assign n8463 = n8408 ^ n8368 ;
  assign n7069 = n6982 ^ n6942 ;
  assign n8464 = n8463 ^ n7069 ;
  assign n4036 = n4031 ^ n4029 ;
  assign n4037 = n4032 ^ n4030 ;
  assign n4038 = n4036 & n4037 ;
  assign n4040 = n4038 ^ n4034 ;
  assign n4045 = n4042 ^ n4040 ;
  assign n4033 = n4028 ^ n4027 ;
  assign n4046 = n4045 ^ n4033 ;
  assign n4057 = n4050 ^ n4046 ;
  assign n4012 = n4003 ^ n4001 ;
  assign n4014 = n4012 ^ n3999 ;
  assign n4058 = n4057 ^ n4014 ;
  assign n3917 = n3912 ^ n3910 ;
  assign n3918 = n3913 ^ n3911 ;
  assign n3919 = n3917 & n3918 ;
  assign n3921 = n3919 ^ n3915 ;
  assign n3926 = n3923 ^ n3921 ;
  assign n3914 = n3909 ^ n3908 ;
  assign n3927 = n3926 ^ n3914 ;
  assign n3938 = n3931 ^ n3927 ;
  assign n3893 = n3884 ^ n3882 ;
  assign n3895 = n3893 ^ n3880 ;
  assign n3939 = n3938 ^ n3895 ;
  assign n4208 = n4058 ^ n3939 ;
  assign n4255 = n4232 ^ n4208 ;
  assign n4256 = n4255 ^ n3773 ;
  assign n4351 = n4296 ^ n4256 ;
  assign n2957 = n2870 ^ n2830 ;
  assign n4352 = n4351 ^ n2957 ;
  assign n12839 = n8464 ^ n4352 ;
  assign n8185 = n7916 ^ n7900 ;
  assign n8186 = n7917 ^ n7901 ;
  assign n8234 = n8185 & n8186 ;
  assign n8183 = n7914 ^ n7898 ;
  assign n8184 = n7915 ^ n7899 ;
  assign n8233 = n8183 & n8184 ;
  assign n8238 = n8234 ^ n8233 ;
  assign n8181 = n7912 ^ n7896 ;
  assign n8182 = n7913 ^ n7897 ;
  assign n8227 = n8181 & n8182 ;
  assign n8179 = n7910 ^ n7894 ;
  assign n8180 = n7911 ^ n7895 ;
  assign n8226 = n8179 & n8180 ;
  assign n8231 = n8227 ^ n8226 ;
  assign n8252 = n8238 ^ n8231 ;
  assign n8177 = n7908 ^ n7892 ;
  assign n8178 = n7909 ^ n7893 ;
  assign n8202 = n8177 & n8178 ;
  assign n8175 = n7906 ^ n7890 ;
  assign n8176 = n7907 ^ n7891 ;
  assign n8201 = n8175 & n8176 ;
  assign n8206 = n8202 ^ n8201 ;
  assign n8173 = n7904 ^ n7888 ;
  assign n8174 = n7905 ^ n7889 ;
  assign n8195 = n8173 & n8174 ;
  assign n8171 = n7902 ^ n7886 ;
  assign n8172 = n7903 ^ n7887 ;
  assign n8194 = n8171 & n8172 ;
  assign n8199 = n8195 ^ n8194 ;
  assign n8220 = n8206 ^ n8199 ;
  assign n8301 = n8252 ^ n8220 ;
  assign n8321 = n8313 ^ n8301 ;
  assign n8322 = n8321 ^ n8164 ;
  assign n8369 = n8345 ^ n8322 ;
  assign n7925 = n7879 ^ n7862 ;
  assign n8370 = n8369 ^ n7925 ;
  assign n8465 = n8409 ^ n8370 ;
  assign n7054 = n6976 ^ n6952 ;
  assign n7070 = n7054 ^ n6943 ;
  assign n8466 = n8465 ^ n7070 ;
  assign n4073 = n3804 ^ n3788 ;
  assign n4074 = n3805 ^ n3789 ;
  assign n4122 = n4073 & n4074 ;
  assign n4071 = n3802 ^ n3786 ;
  assign n4072 = n3803 ^ n3787 ;
  assign n4121 = n4071 & n4072 ;
  assign n4126 = n4122 ^ n4121 ;
  assign n4069 = n3800 ^ n3784 ;
  assign n4070 = n3801 ^ n3785 ;
  assign n4115 = n4069 & n4070 ;
  assign n4067 = n3798 ^ n3782 ;
  assign n4068 = n3799 ^ n3783 ;
  assign n4114 = n4067 & n4068 ;
  assign n4119 = n4115 ^ n4114 ;
  assign n4140 = n4126 ^ n4119 ;
  assign n4065 = n3796 ^ n3780 ;
  assign n4066 = n3797 ^ n3781 ;
  assign n4090 = n4065 & n4066 ;
  assign n4063 = n3794 ^ n3778 ;
  assign n4064 = n3795 ^ n3779 ;
  assign n4089 = n4063 & n4064 ;
  assign n4094 = n4090 ^ n4089 ;
  assign n4061 = n3792 ^ n3776 ;
  assign n4062 = n3793 ^ n3777 ;
  assign n4083 = n4061 & n4062 ;
  assign n4059 = n3790 ^ n3774 ;
  assign n4060 = n3791 ^ n3775 ;
  assign n4082 = n4059 & n4060 ;
  assign n4087 = n4083 ^ n4082 ;
  assign n4108 = n4094 ^ n4087 ;
  assign n4189 = n4140 ^ n4108 ;
  assign n4209 = n4201 ^ n4189 ;
  assign n4210 = n4209 ^ n4052 ;
  assign n4257 = n4233 ^ n4210 ;
  assign n3813 = n3767 ^ n3750 ;
  assign n4258 = n4257 ^ n3813 ;
  assign n4353 = n4297 ^ n4258 ;
  assign n2942 = n2864 ^ n2840 ;
  assign n2958 = n2942 ^ n2831 ;
  assign n4354 = n4353 ^ n2958 ;
  assign n12840 = n8466 ^ n4354 ;
  assign n8235 = n8185 ^ n8183 ;
  assign n8236 = n8186 ^ n8184 ;
  assign n8237 = n8235 & n8236 ;
  assign n8239 = n8237 ^ n8233 ;
  assign n8228 = n8181 ^ n8179 ;
  assign n8229 = n8182 ^ n8180 ;
  assign n8230 = n8228 & n8229 ;
  assign n8232 = n8230 ^ n8226 ;
  assign n8253 = n8239 ^ n8232 ;
  assign n8203 = n8177 ^ n8175 ;
  assign n8204 = n8178 ^ n8176 ;
  assign n8205 = n8203 & n8204 ;
  assign n8207 = n8205 ^ n8201 ;
  assign n8196 = n8173 ^ n8171 ;
  assign n8197 = n8174 ^ n8172 ;
  assign n8198 = n8196 & n8197 ;
  assign n8200 = n8198 ^ n8194 ;
  assign n8221 = n8207 ^ n8200 ;
  assign n8302 = n8253 ^ n8221 ;
  assign n8323 = n8314 ^ n8302 ;
  assign n8324 = n8323 ^ n8166 ;
  assign n8371 = n8346 ^ n8324 ;
  assign n7926 = n7881 ^ n7863 ;
  assign n8372 = n8371 ^ n7926 ;
  assign n8467 = n8410 ^ n8372 ;
  assign n7055 = n6978 ^ n6954 ;
  assign n7071 = n7055 ^ n6944 ;
  assign n8468 = n8467 ^ n7071 ;
  assign n4123 = n4073 ^ n4071 ;
  assign n4124 = n4074 ^ n4072 ;
  assign n4125 = n4123 & n4124 ;
  assign n4127 = n4125 ^ n4121 ;
  assign n4116 = n4069 ^ n4067 ;
  assign n4117 = n4070 ^ n4068 ;
  assign n4118 = n4116 & n4117 ;
  assign n4120 = n4118 ^ n4114 ;
  assign n4141 = n4127 ^ n4120 ;
  assign n4091 = n4065 ^ n4063 ;
  assign n4092 = n4066 ^ n4064 ;
  assign n4093 = n4091 & n4092 ;
  assign n4095 = n4093 ^ n4089 ;
  assign n4084 = n4061 ^ n4059 ;
  assign n4085 = n4062 ^ n4060 ;
  assign n4086 = n4084 & n4085 ;
  assign n4088 = n4086 ^ n4082 ;
  assign n4109 = n4095 ^ n4088 ;
  assign n4190 = n4141 ^ n4109 ;
  assign n4211 = n4202 ^ n4190 ;
  assign n4212 = n4211 ^ n4054 ;
  assign n4259 = n4234 ^ n4212 ;
  assign n3814 = n3769 ^ n3751 ;
  assign n4260 = n4259 ^ n3814 ;
  assign n4355 = n4298 ^ n4260 ;
  assign n2943 = n2866 ^ n2842 ;
  assign n2959 = n2943 ^ n2832 ;
  assign n4356 = n4355 ^ n2959 ;
  assign n12841 = n8468 ^ n4356 ;
  assign n8242 = n8185 ^ n8181 ;
  assign n8243 = n8186 ^ n8182 ;
  assign n8246 = n8242 & n8243 ;
  assign n8240 = n8183 ^ n8179 ;
  assign n8241 = n8184 ^ n8180 ;
  assign n8245 = n8240 & n8241 ;
  assign n8250 = n8246 ^ n8245 ;
  assign n8254 = n8252 ^ n8250 ;
  assign n8255 = n8254 ^ n8239 ;
  assign n8210 = n8177 ^ n8173 ;
  assign n8211 = n8178 ^ n8174 ;
  assign n8214 = n8210 & n8211 ;
  assign n8208 = n8175 ^ n8171 ;
  assign n8209 = n8176 ^ n8172 ;
  assign n8213 = n8208 & n8209 ;
  assign n8218 = n8214 ^ n8213 ;
  assign n8222 = n8220 ^ n8218 ;
  assign n8223 = n8222 ^ n8207 ;
  assign n8303 = n8255 ^ n8223 ;
  assign n8325 = n8315 ^ n8303 ;
  assign n8326 = n8325 ^ n8168 ;
  assign n8373 = n8347 ^ n8326 ;
  assign n7927 = n7883 ^ n7864 ;
  assign n8374 = n8373 ^ n7927 ;
  assign n8469 = n8411 ^ n8374 ;
  assign n7056 = n6980 ^ n6956 ;
  assign n7072 = n7056 ^ n6945 ;
  assign n8470 = n8469 ^ n7072 ;
  assign n4130 = n4073 ^ n4069 ;
  assign n4131 = n4074 ^ n4070 ;
  assign n4134 = n4130 & n4131 ;
  assign n4128 = n4071 ^ n4067 ;
  assign n4129 = n4072 ^ n4068 ;
  assign n4133 = n4128 & n4129 ;
  assign n4138 = n4134 ^ n4133 ;
  assign n4142 = n4140 ^ n4138 ;
  assign n4143 = n4142 ^ n4127 ;
  assign n4098 = n4065 ^ n4061 ;
  assign n4099 = n4066 ^ n4062 ;
  assign n4102 = n4098 & n4099 ;
  assign n4096 = n4063 ^ n4059 ;
  assign n4097 = n4064 ^ n4060 ;
  assign n4101 = n4096 & n4097 ;
  assign n4106 = n4102 ^ n4101 ;
  assign n4110 = n4108 ^ n4106 ;
  assign n4111 = n4110 ^ n4095 ;
  assign n4191 = n4143 ^ n4111 ;
  assign n4213 = n4203 ^ n4191 ;
  assign n4214 = n4213 ^ n4056 ;
  assign n4261 = n4235 ^ n4214 ;
  assign n3815 = n3771 ^ n3752 ;
  assign n4262 = n4261 ^ n3815 ;
  assign n4357 = n4299 ^ n4262 ;
  assign n2944 = n2868 ^ n2844 ;
  assign n2960 = n2944 ^ n2833 ;
  assign n4358 = n4357 ^ n2960 ;
  assign n12842 = n8470 ^ n4358 ;
  assign n8247 = n8242 ^ n8240 ;
  assign n8248 = n8243 ^ n8241 ;
  assign n8249 = n8247 & n8248 ;
  assign n8251 = n8249 ^ n8245 ;
  assign n8256 = n8253 ^ n8251 ;
  assign n8244 = n8239 ^ n8238 ;
  assign n8257 = n8256 ^ n8244 ;
  assign n8215 = n8210 ^ n8208 ;
  assign n8216 = n8211 ^ n8209 ;
  assign n8217 = n8215 & n8216 ;
  assign n8219 = n8217 ^ n8213 ;
  assign n8224 = n8221 ^ n8219 ;
  assign n8212 = n8207 ^ n8206 ;
  assign n8225 = n8224 ^ n8212 ;
  assign n8304 = n8257 ^ n8225 ;
  assign n8327 = n8316 ^ n8304 ;
  assign n8328 = n8327 ^ n8170 ;
  assign n8375 = n8348 ^ n8328 ;
  assign n7928 = n7885 ^ n7865 ;
  assign n8376 = n8375 ^ n7928 ;
  assign n8471 = n8412 ^ n8376 ;
  assign n7057 = n6982 ^ n6958 ;
  assign n7073 = n7057 ^ n6946 ;
  assign n8472 = n8471 ^ n7073 ;
  assign n4135 = n4130 ^ n4128 ;
  assign n4136 = n4131 ^ n4129 ;
  assign n4137 = n4135 & n4136 ;
  assign n4139 = n4137 ^ n4133 ;
  assign n4144 = n4141 ^ n4139 ;
  assign n4132 = n4127 ^ n4126 ;
  assign n4145 = n4144 ^ n4132 ;
  assign n4103 = n4098 ^ n4096 ;
  assign n4104 = n4099 ^ n4097 ;
  assign n4105 = n4103 & n4104 ;
  assign n4107 = n4105 ^ n4101 ;
  assign n4112 = n4109 ^ n4107 ;
  assign n4100 = n4095 ^ n4094 ;
  assign n4113 = n4112 ^ n4100 ;
  assign n4192 = n4145 ^ n4113 ;
  assign n4215 = n4204 ^ n4192 ;
  assign n4216 = n4215 ^ n4058 ;
  assign n4263 = n4236 ^ n4216 ;
  assign n3816 = n3773 ^ n3753 ;
  assign n4264 = n4263 ^ n3816 ;
  assign n4359 = n4300 ^ n4264 ;
  assign n2945 = n2870 ^ n2846 ;
  assign n2961 = n2945 ^ n2834 ;
  assign n4360 = n4359 ^ n2961 ;
  assign n12843 = n8472 ^ n4360 ;
  assign n8264 = n8185 ^ n8177 ;
  assign n8265 = n8186 ^ n8178 ;
  assign n8277 = n8264 & n8265 ;
  assign n8262 = n8183 ^ n8175 ;
  assign n8263 = n8184 ^ n8176 ;
  assign n8276 = n8262 & n8263 ;
  assign n8281 = n8277 ^ n8276 ;
  assign n8260 = n8181 ^ n8173 ;
  assign n8261 = n8182 ^ n8174 ;
  assign n8270 = n8260 & n8261 ;
  assign n8258 = n8179 ^ n8171 ;
  assign n8259 = n8180 ^ n8172 ;
  assign n8269 = n8258 & n8259 ;
  assign n8274 = n8270 ^ n8269 ;
  assign n8295 = n8281 ^ n8274 ;
  assign n8305 = n8301 ^ n8295 ;
  assign n8306 = n8305 ^ n8255 ;
  assign n8329 = n8317 ^ n8306 ;
  assign n8190 = n8168 ^ n8159 ;
  assign n8330 = n8329 ^ n8190 ;
  assign n8377 = n8349 ^ n8330 ;
  assign n7921 = n7883 ^ n7871 ;
  assign n7929 = n7921 ^ n7866 ;
  assign n8378 = n8377 ^ n7929 ;
  assign n8473 = n8413 ^ n8378 ;
  assign n7050 = n6980 ^ n6968 ;
  assign n7058 = n7050 ^ n6960 ;
  assign n7074 = n7058 ^ n6947 ;
  assign n8474 = n8473 ^ n7074 ;
  assign n4152 = n4073 ^ n4065 ;
  assign n4153 = n4074 ^ n4066 ;
  assign n4165 = n4152 & n4153 ;
  assign n4150 = n4071 ^ n4063 ;
  assign n4151 = n4072 ^ n4064 ;
  assign n4164 = n4150 & n4151 ;
  assign n4169 = n4165 ^ n4164 ;
  assign n4148 = n4069 ^ n4061 ;
  assign n4149 = n4070 ^ n4062 ;
  assign n4158 = n4148 & n4149 ;
  assign n4146 = n4067 ^ n4059 ;
  assign n4147 = n4068 ^ n4060 ;
  assign n4157 = n4146 & n4147 ;
  assign n4162 = n4158 ^ n4157 ;
  assign n4183 = n4169 ^ n4162 ;
  assign n4193 = n4189 ^ n4183 ;
  assign n4194 = n4193 ^ n4143 ;
  assign n4217 = n4205 ^ n4194 ;
  assign n4078 = n4056 ^ n4047 ;
  assign n4218 = n4217 ^ n4078 ;
  assign n4265 = n4237 ^ n4218 ;
  assign n3809 = n3771 ^ n3759 ;
  assign n3817 = n3809 ^ n3754 ;
  assign n4266 = n4265 ^ n3817 ;
  assign n4361 = n4301 ^ n4266 ;
  assign n2938 = n2868 ^ n2856 ;
  assign n2946 = n2938 ^ n2848 ;
  assign n2962 = n2946 ^ n2835 ;
  assign n4362 = n4361 ^ n2962 ;
  assign n12844 = n8474 ^ n4362 ;
  assign n8278 = n8264 ^ n8262 ;
  assign n8279 = n8265 ^ n8263 ;
  assign n8280 = n8278 & n8279 ;
  assign n8282 = n8280 ^ n8276 ;
  assign n8271 = n8260 ^ n8258 ;
  assign n8272 = n8261 ^ n8259 ;
  assign n8273 = n8271 & n8272 ;
  assign n8275 = n8273 ^ n8269 ;
  assign n8296 = n8282 ^ n8275 ;
  assign n8307 = n8302 ^ n8296 ;
  assign n8308 = n8307 ^ n8257 ;
  assign n8331 = n8318 ^ n8308 ;
  assign n8191 = n8170 ^ n8160 ;
  assign n8332 = n8331 ^ n8191 ;
  assign n8379 = n8350 ^ n8332 ;
  assign n7922 = n7885 ^ n7873 ;
  assign n7930 = n7922 ^ n7867 ;
  assign n8380 = n8379 ^ n7930 ;
  assign n8475 = n8414 ^ n8380 ;
  assign n7051 = n6982 ^ n6970 ;
  assign n7059 = n7051 ^ n6962 ;
  assign n7075 = n7059 ^ n6948 ;
  assign n8476 = n8475 ^ n7075 ;
  assign n4166 = n4152 ^ n4150 ;
  assign n4167 = n4153 ^ n4151 ;
  assign n4168 = n4166 & n4167 ;
  assign n4170 = n4168 ^ n4164 ;
  assign n4159 = n4148 ^ n4146 ;
  assign n4160 = n4149 ^ n4147 ;
  assign n4161 = n4159 & n4160 ;
  assign n4163 = n4161 ^ n4157 ;
  assign n4184 = n4170 ^ n4163 ;
  assign n4195 = n4190 ^ n4184 ;
  assign n4196 = n4195 ^ n4145 ;
  assign n4219 = n4206 ^ n4196 ;
  assign n4079 = n4058 ^ n4048 ;
  assign n4220 = n4219 ^ n4079 ;
  assign n4267 = n4238 ^ n4220 ;
  assign n3810 = n3773 ^ n3761 ;
  assign n3818 = n3810 ^ n3755 ;
  assign n4268 = n4267 ^ n3818 ;
  assign n4363 = n4302 ^ n4268 ;
  assign n2939 = n2870 ^ n2858 ;
  assign n2947 = n2939 ^ n2850 ;
  assign n2963 = n2947 ^ n2836 ;
  assign n4364 = n4363 ^ n2963 ;
  assign n12845 = n8476 ^ n4364 ;
  assign n8285 = n8264 ^ n8260 ;
  assign n8286 = n8265 ^ n8261 ;
  assign n8289 = n8285 & n8286 ;
  assign n8283 = n8262 ^ n8258 ;
  assign n8284 = n8263 ^ n8259 ;
  assign n8288 = n8283 & n8284 ;
  assign n8293 = n8289 ^ n8288 ;
  assign n8297 = n8295 ^ n8293 ;
  assign n8298 = n8297 ^ n8282 ;
  assign n8309 = n8303 ^ n8298 ;
  assign n8267 = n8257 ^ n8252 ;
  assign n8310 = n8309 ^ n8267 ;
  assign n8333 = n8319 ^ n8310 ;
  assign n8188 = n8170 ^ n8164 ;
  assign n8192 = n8188 ^ n8161 ;
  assign n8334 = n8333 ^ n8192 ;
  assign n8381 = n8351 ^ n8334 ;
  assign n7919 = n7885 ^ n7879 ;
  assign n7923 = n7919 ^ n7875 ;
  assign n7931 = n7923 ^ n7868 ;
  assign n8382 = n8381 ^ n7931 ;
  assign n8477 = n8415 ^ n8382 ;
  assign n7048 = n6982 ^ n6976 ;
  assign n7052 = n7048 ^ n6972 ;
  assign n7060 = n7052 ^ n6964 ;
  assign n7076 = n7060 ^ n6949 ;
  assign n8478 = n8477 ^ n7076 ;
  assign n4173 = n4152 ^ n4148 ;
  assign n4174 = n4153 ^ n4149 ;
  assign n4177 = n4173 & n4174 ;
  assign n4171 = n4150 ^ n4146 ;
  assign n4172 = n4151 ^ n4147 ;
  assign n4176 = n4171 & n4172 ;
  assign n4181 = n4177 ^ n4176 ;
  assign n4185 = n4183 ^ n4181 ;
  assign n4186 = n4185 ^ n4170 ;
  assign n4197 = n4191 ^ n4186 ;
  assign n4155 = n4145 ^ n4140 ;
  assign n4198 = n4197 ^ n4155 ;
  assign n4221 = n4207 ^ n4198 ;
  assign n4076 = n4058 ^ n4052 ;
  assign n4080 = n4076 ^ n4049 ;
  assign n4222 = n4221 ^ n4080 ;
  assign n4269 = n4239 ^ n4222 ;
  assign n3807 = n3773 ^ n3767 ;
  assign n3811 = n3807 ^ n3763 ;
  assign n3819 = n3811 ^ n3756 ;
  assign n4270 = n4269 ^ n3819 ;
  assign n4365 = n4303 ^ n4270 ;
  assign n2936 = n2870 ^ n2864 ;
  assign n2940 = n2936 ^ n2860 ;
  assign n2948 = n2940 ^ n2852 ;
  assign n2964 = n2948 ^ n2837 ;
  assign n4366 = n4365 ^ n2964 ;
  assign n12846 = n8478 ^ n4366 ;
  assign n8290 = n8285 ^ n8283 ;
  assign n8291 = n8286 ^ n8284 ;
  assign n8292 = n8290 & n8291 ;
  assign n8294 = n8292 ^ n8288 ;
  assign n8299 = n8296 ^ n8294 ;
  assign n8287 = n8282 ^ n8281 ;
  assign n8300 = n8299 ^ n8287 ;
  assign n8311 = n8304 ^ n8300 ;
  assign n8266 = n8257 ^ n8255 ;
  assign n8268 = n8266 ^ n8253 ;
  assign n8312 = n8311 ^ n8268 ;
  assign n8335 = n8320 ^ n8312 ;
  assign n8187 = n8170 ^ n8168 ;
  assign n8189 = n8187 ^ n8166 ;
  assign n8193 = n8189 ^ n8162 ;
  assign n8336 = n8335 ^ n8193 ;
  assign n8383 = n8352 ^ n8336 ;
  assign n7918 = n7885 ^ n7883 ;
  assign n7920 = n7918 ^ n7881 ;
  assign n7924 = n7920 ^ n7877 ;
  assign n7932 = n7924 ^ n7869 ;
  assign n8384 = n8383 ^ n7932 ;
  assign n8479 = n8416 ^ n8384 ;
  assign n7047 = n6982 ^ n6980 ;
  assign n7049 = n7047 ^ n6978 ;
  assign n7053 = n7049 ^ n6974 ;
  assign n7061 = n7053 ^ n6966 ;
  assign n7077 = n7061 ^ n6950 ;
  assign n8480 = n8479 ^ n7077 ;
  assign n4178 = n4173 ^ n4171 ;
  assign n4179 = n4174 ^ n4172 ;
  assign n4180 = n4178 & n4179 ;
  assign n4182 = n4180 ^ n4176 ;
  assign n4187 = n4184 ^ n4182 ;
  assign n4175 = n4170 ^ n4169 ;
  assign n4188 = n4187 ^ n4175 ;
  assign n4199 = n4192 ^ n4188 ;
  assign n4154 = n4145 ^ n4143 ;
  assign n4156 = n4154 ^ n4141 ;
  assign n4200 = n4199 ^ n4156 ;
  assign n4223 = n4208 ^ n4200 ;
  assign n4075 = n4058 ^ n4056 ;
  assign n4077 = n4075 ^ n4054 ;
  assign n4081 = n4077 ^ n4050 ;
  assign n4224 = n4223 ^ n4081 ;
  assign n4271 = n4240 ^ n4224 ;
  assign n3806 = n3773 ^ n3771 ;
  assign n3808 = n3806 ^ n3769 ;
  assign n3812 = n3808 ^ n3765 ;
  assign n3820 = n3812 ^ n3757 ;
  assign n4272 = n4271 ^ n3820 ;
  assign n4367 = n4304 ^ n4272 ;
  assign n2935 = n2870 ^ n2868 ;
  assign n2937 = n2935 ^ n2866 ;
  assign n2941 = n2937 ^ n2862 ;
  assign n2949 = n2941 ^ n2854 ;
  assign n2965 = n2949 ^ n2838 ;
  assign n4368 = n4367 ^ n2965 ;
  assign n12847 = n8480 ^ n4368 ;
  assign n8607 = x127 ^ x63 ;
  assign n8608 = x255 ^ x191 ;
  assign n10542 = n8607 & n8608 ;
  assign n8605 = x126 ^ x62 ;
  assign n8606 = x254 ^ x190 ;
  assign n10541 = n8605 & n8606 ;
  assign n10546 = n10542 ^ n10541 ;
  assign n8603 = x125 ^ x61 ;
  assign n8604 = x253 ^ x189 ;
  assign n10535 = n8603 & n8604 ;
  assign n8601 = x124 ^ x60 ;
  assign n8602 = x252 ^ x188 ;
  assign n10534 = n8601 & n8602 ;
  assign n10539 = n10535 ^ n10534 ;
  assign n10560 = n10546 ^ n10539 ;
  assign n8599 = x123 ^ x59 ;
  assign n8600 = x251 ^ x187 ;
  assign n10510 = n8599 & n8600 ;
  assign n8597 = x122 ^ x58 ;
  assign n8598 = x250 ^ x186 ;
  assign n10509 = n8597 & n8598 ;
  assign n10514 = n10510 ^ n10509 ;
  assign n8595 = x121 ^ x57 ;
  assign n8596 = x249 ^ x185 ;
  assign n10503 = n8595 & n8596 ;
  assign n8593 = x120 ^ x56 ;
  assign n8594 = x248 ^ x184 ;
  assign n10502 = n8593 & n8594 ;
  assign n10507 = n10503 ^ n10502 ;
  assign n10528 = n10514 ^ n10507 ;
  assign n10609 = n10560 ^ n10528 ;
  assign n8591 = x119 ^ x55 ;
  assign n8592 = x247 ^ x183 ;
  assign n10423 = n8591 & n8592 ;
  assign n8589 = x118 ^ x54 ;
  assign n8590 = x246 ^ x182 ;
  assign n10422 = n8589 & n8590 ;
  assign n10427 = n10423 ^ n10422 ;
  assign n8587 = x117 ^ x53 ;
  assign n8588 = x245 ^ x181 ;
  assign n10416 = n8587 & n8588 ;
  assign n8585 = x116 ^ x52 ;
  assign n8586 = x244 ^ x180 ;
  assign n10415 = n8585 & n8586 ;
  assign n10420 = n10416 ^ n10415 ;
  assign n10441 = n10427 ^ n10420 ;
  assign n8583 = x115 ^ x51 ;
  assign n8584 = x243 ^ x179 ;
  assign n10391 = n8583 & n8584 ;
  assign n8581 = x114 ^ x50 ;
  assign n8582 = x242 ^ x178 ;
  assign n10390 = n8581 & n8582 ;
  assign n10395 = n10391 ^ n10390 ;
  assign n8579 = x113 ^ x49 ;
  assign n8580 = x241 ^ x177 ;
  assign n10384 = n8579 & n8580 ;
  assign n8577 = x112 ^ x48 ;
  assign n8578 = x240 ^ x176 ;
  assign n10383 = n8577 & n8578 ;
  assign n10388 = n10384 ^ n10383 ;
  assign n10409 = n10395 ^ n10388 ;
  assign n10490 = n10441 ^ n10409 ;
  assign n10763 = n10609 ^ n10490 ;
  assign n8575 = x111 ^ x47 ;
  assign n8576 = x239 ^ x175 ;
  assign n10138 = n8575 & n8576 ;
  assign n8573 = x110 ^ x46 ;
  assign n8574 = x238 ^ x174 ;
  assign n10137 = n8573 & n8574 ;
  assign n10142 = n10138 ^ n10137 ;
  assign n8571 = x109 ^ x45 ;
  assign n8572 = x237 ^ x173 ;
  assign n10131 = n8571 & n8572 ;
  assign n8569 = x108 ^ x44 ;
  assign n8570 = x236 ^ x172 ;
  assign n10130 = n8569 & n8570 ;
  assign n10135 = n10131 ^ n10130 ;
  assign n10156 = n10142 ^ n10135 ;
  assign n8567 = x107 ^ x43 ;
  assign n8568 = x235 ^ x171 ;
  assign n10106 = n8567 & n8568 ;
  assign n8565 = x106 ^ x42 ;
  assign n8566 = x234 ^ x170 ;
  assign n10105 = n8565 & n8566 ;
  assign n10110 = n10106 ^ n10105 ;
  assign n8563 = x105 ^ x41 ;
  assign n8564 = x233 ^ x169 ;
  assign n10099 = n8563 & n8564 ;
  assign n8561 = x104 ^ x40 ;
  assign n8562 = x232 ^ x168 ;
  assign n10098 = n8561 & n8562 ;
  assign n10103 = n10099 ^ n10098 ;
  assign n10124 = n10110 ^ n10103 ;
  assign n10205 = n10156 ^ n10124 ;
  assign n8559 = x103 ^ x39 ;
  assign n8560 = x231 ^ x167 ;
  assign n10019 = n8559 & n8560 ;
  assign n8557 = x102 ^ x38 ;
  assign n8558 = x230 ^ x166 ;
  assign n10018 = n8557 & n8558 ;
  assign n10023 = n10019 ^ n10018 ;
  assign n8555 = x101 ^ x37 ;
  assign n8556 = x229 ^ x165 ;
  assign n10012 = n8555 & n8556 ;
  assign n8553 = x100 ^ x36 ;
  assign n8554 = x228 ^ x164 ;
  assign n10011 = n8553 & n8554 ;
  assign n10016 = n10012 ^ n10011 ;
  assign n10037 = n10023 ^ n10016 ;
  assign n8551 = x99 ^ x35 ;
  assign n8552 = x227 ^ x163 ;
  assign n9987 = n8551 & n8552 ;
  assign n8549 = x98 ^ x34 ;
  assign n8550 = x226 ^ x162 ;
  assign n9986 = n8549 & n8550 ;
  assign n9991 = n9987 ^ n9986 ;
  assign n8547 = x97 ^ x33 ;
  assign n8548 = x225 ^ x161 ;
  assign n9980 = n8547 & n8548 ;
  assign n8545 = x96 ^ x32 ;
  assign n8546 = x224 ^ x160 ;
  assign n9979 = n8545 & n8546 ;
  assign n9984 = n9980 ^ n9979 ;
  assign n10005 = n9991 ^ n9984 ;
  assign n10086 = n10037 ^ n10005 ;
  assign n10359 = n10205 ^ n10086 ;
  assign n11238 = n10763 ^ n10359 ;
  assign n8543 = x95 ^ x31 ;
  assign n8544 = x223 ^ x159 ;
  assign n9235 = n8543 & n8544 ;
  assign n8541 = x94 ^ x30 ;
  assign n8542 = x222 ^ x158 ;
  assign n9234 = n8541 & n8542 ;
  assign n9239 = n9235 ^ n9234 ;
  assign n8539 = x93 ^ x29 ;
  assign n8540 = x221 ^ x157 ;
  assign n9228 = n8539 & n8540 ;
  assign n8537 = x92 ^ x28 ;
  assign n8538 = x220 ^ x156 ;
  assign n9227 = n8537 & n8538 ;
  assign n9232 = n9228 ^ n9227 ;
  assign n9253 = n9239 ^ n9232 ;
  assign n8535 = x91 ^ x27 ;
  assign n8536 = x219 ^ x155 ;
  assign n9203 = n8535 & n8536 ;
  assign n8533 = x90 ^ x26 ;
  assign n8534 = x218 ^ x154 ;
  assign n9202 = n8533 & n8534 ;
  assign n9207 = n9203 ^ n9202 ;
  assign n8531 = x89 ^ x25 ;
  assign n8532 = x217 ^ x153 ;
  assign n9196 = n8531 & n8532 ;
  assign n8529 = x88 ^ x24 ;
  assign n8530 = x216 ^ x152 ;
  assign n9195 = n8529 & n8530 ;
  assign n9200 = n9196 ^ n9195 ;
  assign n9221 = n9207 ^ n9200 ;
  assign n9302 = n9253 ^ n9221 ;
  assign n8527 = x87 ^ x23 ;
  assign n8528 = x215 ^ x151 ;
  assign n9116 = n8527 & n8528 ;
  assign n8525 = x86 ^ x22 ;
  assign n8526 = x214 ^ x150 ;
  assign n9115 = n8525 & n8526 ;
  assign n9120 = n9116 ^ n9115 ;
  assign n8523 = x85 ^ x21 ;
  assign n8524 = x213 ^ x149 ;
  assign n9109 = n8523 & n8524 ;
  assign n8521 = x84 ^ x20 ;
  assign n8522 = x212 ^ x148 ;
  assign n9108 = n8521 & n8522 ;
  assign n9113 = n9109 ^ n9108 ;
  assign n9134 = n9120 ^ n9113 ;
  assign n8519 = x83 ^ x19 ;
  assign n8520 = x211 ^ x147 ;
  assign n9084 = n8519 & n8520 ;
  assign n8517 = x82 ^ x18 ;
  assign n8518 = x210 ^ x146 ;
  assign n9083 = n8517 & n8518 ;
  assign n9088 = n9084 ^ n9083 ;
  assign n8515 = x81 ^ x17 ;
  assign n8516 = x209 ^ x145 ;
  assign n9077 = n8515 & n8516 ;
  assign n8513 = x80 ^ x16 ;
  assign n8514 = x208 ^ x144 ;
  assign n9076 = n8513 & n8514 ;
  assign n9081 = n9077 ^ n9076 ;
  assign n9102 = n9088 ^ n9081 ;
  assign n9183 = n9134 ^ n9102 ;
  assign n9456 = n9302 ^ n9183 ;
  assign n8511 = x79 ^ x15 ;
  assign n8512 = x207 ^ x143 ;
  assign n8831 = n8511 & n8512 ;
  assign n8509 = x78 ^ x14 ;
  assign n8510 = x206 ^ x142 ;
  assign n8830 = n8509 & n8510 ;
  assign n8835 = n8831 ^ n8830 ;
  assign n8507 = x77 ^ x13 ;
  assign n8508 = x205 ^ x141 ;
  assign n8824 = n8507 & n8508 ;
  assign n8505 = x76 ^ x12 ;
  assign n8506 = x204 ^ x140 ;
  assign n8823 = n8505 & n8506 ;
  assign n8828 = n8824 ^ n8823 ;
  assign n8849 = n8835 ^ n8828 ;
  assign n8503 = x75 ^ x11 ;
  assign n8504 = x203 ^ x139 ;
  assign n8799 = n8503 & n8504 ;
  assign n8501 = x74 ^ x10 ;
  assign n8502 = x202 ^ x138 ;
  assign n8798 = n8501 & n8502 ;
  assign n8803 = n8799 ^ n8798 ;
  assign n8499 = x73 ^ x9 ;
  assign n8500 = x201 ^ x137 ;
  assign n8792 = n8499 & n8500 ;
  assign n8497 = x72 ^ x8 ;
  assign n8498 = x200 ^ x136 ;
  assign n8791 = n8497 & n8498 ;
  assign n8796 = n8792 ^ n8791 ;
  assign n8817 = n8803 ^ n8796 ;
  assign n8898 = n8849 ^ n8817 ;
  assign n8495 = x71 ^ x7 ;
  assign n8496 = x199 ^ x135 ;
  assign n8712 = n8495 & n8496 ;
  assign n8493 = x70 ^ x6 ;
  assign n8494 = x198 ^ x134 ;
  assign n8711 = n8493 & n8494 ;
  assign n8716 = n8712 ^ n8711 ;
  assign n8491 = x69 ^ x5 ;
  assign n8492 = x197 ^ x133 ;
  assign n8705 = n8491 & n8492 ;
  assign n8489 = x68 ^ x4 ;
  assign n8490 = x196 ^ x132 ;
  assign n8704 = n8489 & n8490 ;
  assign n8709 = n8705 ^ n8704 ;
  assign n8730 = n8716 ^ n8709 ;
  assign n8487 = x67 ^ x3 ;
  assign n8488 = x195 ^ x131 ;
  assign n8680 = n8487 & n8488 ;
  assign n8485 = x66 ^ x2 ;
  assign n8486 = x194 ^ x130 ;
  assign n8679 = n8485 & n8486 ;
  assign n8684 = n8680 ^ n8679 ;
  assign n8483 = x65 ^ x1 ;
  assign n8484 = x193 ^ x129 ;
  assign n8673 = n8483 & n8484 ;
  assign n8481 = x64 ^ x0 ;
  assign n8482 = x192 ^ x128 ;
  assign n8672 = n8481 & n8482 ;
  assign n8677 = n8673 ^ n8672 ;
  assign n8698 = n8684 ^ n8677 ;
  assign n8779 = n8730 ^ n8698 ;
  assign n9052 = n8898 ^ n8779 ;
  assign n9931 = n9456 ^ n9052 ;
  assign n12688 = n11238 ^ n9931 ;
  assign n12848 = n12784 ^ n12688 ;
  assign n12849 = n12848 ^ n8418 ;
  assign n10543 = n8607 ^ n8605 ;
  assign n10544 = n8608 ^ n8606 ;
  assign n10545 = n10543 & n10544 ;
  assign n10547 = n10545 ^ n10541 ;
  assign n10536 = n8603 ^ n8601 ;
  assign n10537 = n8604 ^ n8602 ;
  assign n10538 = n10536 & n10537 ;
  assign n10540 = n10538 ^ n10534 ;
  assign n10561 = n10547 ^ n10540 ;
  assign n10511 = n8599 ^ n8597 ;
  assign n10512 = n8600 ^ n8598 ;
  assign n10513 = n10511 & n10512 ;
  assign n10515 = n10513 ^ n10509 ;
  assign n10504 = n8595 ^ n8593 ;
  assign n10505 = n8596 ^ n8594 ;
  assign n10506 = n10504 & n10505 ;
  assign n10508 = n10506 ^ n10502 ;
  assign n10529 = n10515 ^ n10508 ;
  assign n10610 = n10561 ^ n10529 ;
  assign n10424 = n8591 ^ n8589 ;
  assign n10425 = n8592 ^ n8590 ;
  assign n10426 = n10424 & n10425 ;
  assign n10428 = n10426 ^ n10422 ;
  assign n10417 = n8587 ^ n8585 ;
  assign n10418 = n8588 ^ n8586 ;
  assign n10419 = n10417 & n10418 ;
  assign n10421 = n10419 ^ n10415 ;
  assign n10442 = n10428 ^ n10421 ;
  assign n10392 = n8583 ^ n8581 ;
  assign n10393 = n8584 ^ n8582 ;
  assign n10394 = n10392 & n10393 ;
  assign n10396 = n10394 ^ n10390 ;
  assign n10385 = n8579 ^ n8577 ;
  assign n10386 = n8580 ^ n8578 ;
  assign n10387 = n10385 & n10386 ;
  assign n10389 = n10387 ^ n10383 ;
  assign n10410 = n10396 ^ n10389 ;
  assign n10491 = n10442 ^ n10410 ;
  assign n10764 = n10610 ^ n10491 ;
  assign n10139 = n8575 ^ n8573 ;
  assign n10140 = n8576 ^ n8574 ;
  assign n10141 = n10139 & n10140 ;
  assign n10143 = n10141 ^ n10137 ;
  assign n10132 = n8571 ^ n8569 ;
  assign n10133 = n8572 ^ n8570 ;
  assign n10134 = n10132 & n10133 ;
  assign n10136 = n10134 ^ n10130 ;
  assign n10157 = n10143 ^ n10136 ;
  assign n10107 = n8567 ^ n8565 ;
  assign n10108 = n8568 ^ n8566 ;
  assign n10109 = n10107 & n10108 ;
  assign n10111 = n10109 ^ n10105 ;
  assign n10100 = n8563 ^ n8561 ;
  assign n10101 = n8564 ^ n8562 ;
  assign n10102 = n10100 & n10101 ;
  assign n10104 = n10102 ^ n10098 ;
  assign n10125 = n10111 ^ n10104 ;
  assign n10206 = n10157 ^ n10125 ;
  assign n10020 = n8559 ^ n8557 ;
  assign n10021 = n8560 ^ n8558 ;
  assign n10022 = n10020 & n10021 ;
  assign n10024 = n10022 ^ n10018 ;
  assign n10013 = n8555 ^ n8553 ;
  assign n10014 = n8556 ^ n8554 ;
  assign n10015 = n10013 & n10014 ;
  assign n10017 = n10015 ^ n10011 ;
  assign n10038 = n10024 ^ n10017 ;
  assign n9988 = n8551 ^ n8549 ;
  assign n9989 = n8552 ^ n8550 ;
  assign n9990 = n9988 & n9989 ;
  assign n9992 = n9990 ^ n9986 ;
  assign n9981 = n8547 ^ n8545 ;
  assign n9982 = n8548 ^ n8546 ;
  assign n9983 = n9981 & n9982 ;
  assign n9985 = n9983 ^ n9979 ;
  assign n10006 = n9992 ^ n9985 ;
  assign n10087 = n10038 ^ n10006 ;
  assign n10360 = n10206 ^ n10087 ;
  assign n11239 = n10764 ^ n10360 ;
  assign n9236 = n8543 ^ n8541 ;
  assign n9237 = n8544 ^ n8542 ;
  assign n9238 = n9236 & n9237 ;
  assign n9240 = n9238 ^ n9234 ;
  assign n9229 = n8539 ^ n8537 ;
  assign n9230 = n8540 ^ n8538 ;
  assign n9231 = n9229 & n9230 ;
  assign n9233 = n9231 ^ n9227 ;
  assign n9254 = n9240 ^ n9233 ;
  assign n9204 = n8535 ^ n8533 ;
  assign n9205 = n8536 ^ n8534 ;
  assign n9206 = n9204 & n9205 ;
  assign n9208 = n9206 ^ n9202 ;
  assign n9197 = n8531 ^ n8529 ;
  assign n9198 = n8532 ^ n8530 ;
  assign n9199 = n9197 & n9198 ;
  assign n9201 = n9199 ^ n9195 ;
  assign n9222 = n9208 ^ n9201 ;
  assign n9303 = n9254 ^ n9222 ;
  assign n9117 = n8527 ^ n8525 ;
  assign n9118 = n8528 ^ n8526 ;
  assign n9119 = n9117 & n9118 ;
  assign n9121 = n9119 ^ n9115 ;
  assign n9110 = n8523 ^ n8521 ;
  assign n9111 = n8524 ^ n8522 ;
  assign n9112 = n9110 & n9111 ;
  assign n9114 = n9112 ^ n9108 ;
  assign n9135 = n9121 ^ n9114 ;
  assign n9085 = n8519 ^ n8517 ;
  assign n9086 = n8520 ^ n8518 ;
  assign n9087 = n9085 & n9086 ;
  assign n9089 = n9087 ^ n9083 ;
  assign n9078 = n8515 ^ n8513 ;
  assign n9079 = n8516 ^ n8514 ;
  assign n9080 = n9078 & n9079 ;
  assign n9082 = n9080 ^ n9076 ;
  assign n9103 = n9089 ^ n9082 ;
  assign n9184 = n9135 ^ n9103 ;
  assign n9457 = n9303 ^ n9184 ;
  assign n8832 = n8511 ^ n8509 ;
  assign n8833 = n8512 ^ n8510 ;
  assign n8834 = n8832 & n8833 ;
  assign n8836 = n8834 ^ n8830 ;
  assign n8825 = n8507 ^ n8505 ;
  assign n8826 = n8508 ^ n8506 ;
  assign n8827 = n8825 & n8826 ;
  assign n8829 = n8827 ^ n8823 ;
  assign n8850 = n8836 ^ n8829 ;
  assign n8800 = n8503 ^ n8501 ;
  assign n8801 = n8504 ^ n8502 ;
  assign n8802 = n8800 & n8801 ;
  assign n8804 = n8802 ^ n8798 ;
  assign n8793 = n8499 ^ n8497 ;
  assign n8794 = n8500 ^ n8498 ;
  assign n8795 = n8793 & n8794 ;
  assign n8797 = n8795 ^ n8791 ;
  assign n8818 = n8804 ^ n8797 ;
  assign n8899 = n8850 ^ n8818 ;
  assign n8713 = n8495 ^ n8493 ;
  assign n8714 = n8496 ^ n8494 ;
  assign n8715 = n8713 & n8714 ;
  assign n8717 = n8715 ^ n8711 ;
  assign n8706 = n8491 ^ n8489 ;
  assign n8707 = n8492 ^ n8490 ;
  assign n8708 = n8706 & n8707 ;
  assign n8710 = n8708 ^ n8704 ;
  assign n8731 = n8717 ^ n8710 ;
  assign n8681 = n8487 ^ n8485 ;
  assign n8682 = n8488 ^ n8486 ;
  assign n8683 = n8681 & n8682 ;
  assign n8685 = n8683 ^ n8679 ;
  assign n8674 = n8483 ^ n8481 ;
  assign n8675 = n8484 ^ n8482 ;
  assign n8676 = n8674 & n8675 ;
  assign n8678 = n8676 ^ n8672 ;
  assign n8699 = n8685 ^ n8678 ;
  assign n8780 = n8731 ^ n8699 ;
  assign n9053 = n8899 ^ n8780 ;
  assign n9932 = n9457 ^ n9053 ;
  assign n12689 = n11239 ^ n9932 ;
  assign n12850 = n12785 ^ n12689 ;
  assign n12851 = n12850 ^ n8420 ;
  assign n10550 = n8607 ^ n8603 ;
  assign n10551 = n8608 ^ n8604 ;
  assign n10554 = n10550 & n10551 ;
  assign n10548 = n8605 ^ n8601 ;
  assign n10549 = n8606 ^ n8602 ;
  assign n10553 = n10548 & n10549 ;
  assign n10558 = n10554 ^ n10553 ;
  assign n10562 = n10560 ^ n10558 ;
  assign n10563 = n10562 ^ n10547 ;
  assign n10518 = n8599 ^ n8595 ;
  assign n10519 = n8600 ^ n8596 ;
  assign n10522 = n10518 & n10519 ;
  assign n10516 = n8597 ^ n8593 ;
  assign n10517 = n8598 ^ n8594 ;
  assign n10521 = n10516 & n10517 ;
  assign n10526 = n10522 ^ n10521 ;
  assign n10530 = n10528 ^ n10526 ;
  assign n10531 = n10530 ^ n10515 ;
  assign n10611 = n10563 ^ n10531 ;
  assign n10431 = n8591 ^ n8587 ;
  assign n10432 = n8592 ^ n8588 ;
  assign n10435 = n10431 & n10432 ;
  assign n10429 = n8589 ^ n8585 ;
  assign n10430 = n8590 ^ n8586 ;
  assign n10434 = n10429 & n10430 ;
  assign n10439 = n10435 ^ n10434 ;
  assign n10443 = n10441 ^ n10439 ;
  assign n10444 = n10443 ^ n10428 ;
  assign n10399 = n8583 ^ n8579 ;
  assign n10400 = n8584 ^ n8580 ;
  assign n10403 = n10399 & n10400 ;
  assign n10397 = n8581 ^ n8577 ;
  assign n10398 = n8582 ^ n8578 ;
  assign n10402 = n10397 & n10398 ;
  assign n10407 = n10403 ^ n10402 ;
  assign n10411 = n10409 ^ n10407 ;
  assign n10412 = n10411 ^ n10396 ;
  assign n10492 = n10444 ^ n10412 ;
  assign n10765 = n10611 ^ n10492 ;
  assign n10146 = n8575 ^ n8571 ;
  assign n10147 = n8576 ^ n8572 ;
  assign n10150 = n10146 & n10147 ;
  assign n10144 = n8573 ^ n8569 ;
  assign n10145 = n8574 ^ n8570 ;
  assign n10149 = n10144 & n10145 ;
  assign n10154 = n10150 ^ n10149 ;
  assign n10158 = n10156 ^ n10154 ;
  assign n10159 = n10158 ^ n10143 ;
  assign n10114 = n8567 ^ n8563 ;
  assign n10115 = n8568 ^ n8564 ;
  assign n10118 = n10114 & n10115 ;
  assign n10112 = n8565 ^ n8561 ;
  assign n10113 = n8566 ^ n8562 ;
  assign n10117 = n10112 & n10113 ;
  assign n10122 = n10118 ^ n10117 ;
  assign n10126 = n10124 ^ n10122 ;
  assign n10127 = n10126 ^ n10111 ;
  assign n10207 = n10159 ^ n10127 ;
  assign n10027 = n8559 ^ n8555 ;
  assign n10028 = n8560 ^ n8556 ;
  assign n10031 = n10027 & n10028 ;
  assign n10025 = n8557 ^ n8553 ;
  assign n10026 = n8558 ^ n8554 ;
  assign n10030 = n10025 & n10026 ;
  assign n10035 = n10031 ^ n10030 ;
  assign n10039 = n10037 ^ n10035 ;
  assign n10040 = n10039 ^ n10024 ;
  assign n9995 = n8551 ^ n8547 ;
  assign n9996 = n8552 ^ n8548 ;
  assign n9999 = n9995 & n9996 ;
  assign n9993 = n8549 ^ n8545 ;
  assign n9994 = n8550 ^ n8546 ;
  assign n9998 = n9993 & n9994 ;
  assign n10003 = n9999 ^ n9998 ;
  assign n10007 = n10005 ^ n10003 ;
  assign n10008 = n10007 ^ n9992 ;
  assign n10088 = n10040 ^ n10008 ;
  assign n10361 = n10207 ^ n10088 ;
  assign n11240 = n10765 ^ n10361 ;
  assign n9243 = n8543 ^ n8539 ;
  assign n9244 = n8544 ^ n8540 ;
  assign n9247 = n9243 & n9244 ;
  assign n9241 = n8541 ^ n8537 ;
  assign n9242 = n8542 ^ n8538 ;
  assign n9246 = n9241 & n9242 ;
  assign n9251 = n9247 ^ n9246 ;
  assign n9255 = n9253 ^ n9251 ;
  assign n9256 = n9255 ^ n9240 ;
  assign n9211 = n8535 ^ n8531 ;
  assign n9212 = n8536 ^ n8532 ;
  assign n9215 = n9211 & n9212 ;
  assign n9209 = n8533 ^ n8529 ;
  assign n9210 = n8534 ^ n8530 ;
  assign n9214 = n9209 & n9210 ;
  assign n9219 = n9215 ^ n9214 ;
  assign n9223 = n9221 ^ n9219 ;
  assign n9224 = n9223 ^ n9208 ;
  assign n9304 = n9256 ^ n9224 ;
  assign n9124 = n8527 ^ n8523 ;
  assign n9125 = n8528 ^ n8524 ;
  assign n9128 = n9124 & n9125 ;
  assign n9122 = n8525 ^ n8521 ;
  assign n9123 = n8526 ^ n8522 ;
  assign n9127 = n9122 & n9123 ;
  assign n9132 = n9128 ^ n9127 ;
  assign n9136 = n9134 ^ n9132 ;
  assign n9137 = n9136 ^ n9121 ;
  assign n9092 = n8519 ^ n8515 ;
  assign n9093 = n8520 ^ n8516 ;
  assign n9096 = n9092 & n9093 ;
  assign n9090 = n8517 ^ n8513 ;
  assign n9091 = n8518 ^ n8514 ;
  assign n9095 = n9090 & n9091 ;
  assign n9100 = n9096 ^ n9095 ;
  assign n9104 = n9102 ^ n9100 ;
  assign n9105 = n9104 ^ n9089 ;
  assign n9185 = n9137 ^ n9105 ;
  assign n9458 = n9304 ^ n9185 ;
  assign n8839 = n8511 ^ n8507 ;
  assign n8840 = n8512 ^ n8508 ;
  assign n8843 = n8839 & n8840 ;
  assign n8837 = n8509 ^ n8505 ;
  assign n8838 = n8510 ^ n8506 ;
  assign n8842 = n8837 & n8838 ;
  assign n8847 = n8843 ^ n8842 ;
  assign n8851 = n8849 ^ n8847 ;
  assign n8852 = n8851 ^ n8836 ;
  assign n8807 = n8503 ^ n8499 ;
  assign n8808 = n8504 ^ n8500 ;
  assign n8811 = n8807 & n8808 ;
  assign n8805 = n8501 ^ n8497 ;
  assign n8806 = n8502 ^ n8498 ;
  assign n8810 = n8805 & n8806 ;
  assign n8815 = n8811 ^ n8810 ;
  assign n8819 = n8817 ^ n8815 ;
  assign n8820 = n8819 ^ n8804 ;
  assign n8900 = n8852 ^ n8820 ;
  assign n8720 = n8495 ^ n8491 ;
  assign n8721 = n8496 ^ n8492 ;
  assign n8724 = n8720 & n8721 ;
  assign n8718 = n8493 ^ n8489 ;
  assign n8719 = n8494 ^ n8490 ;
  assign n8723 = n8718 & n8719 ;
  assign n8728 = n8724 ^ n8723 ;
  assign n8732 = n8730 ^ n8728 ;
  assign n8733 = n8732 ^ n8717 ;
  assign n8688 = n8487 ^ n8483 ;
  assign n8689 = n8488 ^ n8484 ;
  assign n8692 = n8688 & n8689 ;
  assign n8686 = n8485 ^ n8481 ;
  assign n8687 = n8486 ^ n8482 ;
  assign n8691 = n8686 & n8687 ;
  assign n8696 = n8692 ^ n8691 ;
  assign n8700 = n8698 ^ n8696 ;
  assign n8701 = n8700 ^ n8685 ;
  assign n8781 = n8733 ^ n8701 ;
  assign n9054 = n8900 ^ n8781 ;
  assign n9933 = n9458 ^ n9054 ;
  assign n12690 = n11240 ^ n9933 ;
  assign n12852 = n12786 ^ n12690 ;
  assign n12853 = n12852 ^ n8422 ;
  assign n10555 = n10550 ^ n10548 ;
  assign n10556 = n10551 ^ n10549 ;
  assign n10557 = n10555 & n10556 ;
  assign n10559 = n10557 ^ n10553 ;
  assign n10564 = n10561 ^ n10559 ;
  assign n10552 = n10547 ^ n10546 ;
  assign n10565 = n10564 ^ n10552 ;
  assign n10523 = n10518 ^ n10516 ;
  assign n10524 = n10519 ^ n10517 ;
  assign n10525 = n10523 & n10524 ;
  assign n10527 = n10525 ^ n10521 ;
  assign n10532 = n10529 ^ n10527 ;
  assign n10520 = n10515 ^ n10514 ;
  assign n10533 = n10532 ^ n10520 ;
  assign n10612 = n10565 ^ n10533 ;
  assign n10436 = n10431 ^ n10429 ;
  assign n10437 = n10432 ^ n10430 ;
  assign n10438 = n10436 & n10437 ;
  assign n10440 = n10438 ^ n10434 ;
  assign n10445 = n10442 ^ n10440 ;
  assign n10433 = n10428 ^ n10427 ;
  assign n10446 = n10445 ^ n10433 ;
  assign n10404 = n10399 ^ n10397 ;
  assign n10405 = n10400 ^ n10398 ;
  assign n10406 = n10404 & n10405 ;
  assign n10408 = n10406 ^ n10402 ;
  assign n10413 = n10410 ^ n10408 ;
  assign n10401 = n10396 ^ n10395 ;
  assign n10414 = n10413 ^ n10401 ;
  assign n10493 = n10446 ^ n10414 ;
  assign n10766 = n10612 ^ n10493 ;
  assign n10151 = n10146 ^ n10144 ;
  assign n10152 = n10147 ^ n10145 ;
  assign n10153 = n10151 & n10152 ;
  assign n10155 = n10153 ^ n10149 ;
  assign n10160 = n10157 ^ n10155 ;
  assign n10148 = n10143 ^ n10142 ;
  assign n10161 = n10160 ^ n10148 ;
  assign n10119 = n10114 ^ n10112 ;
  assign n10120 = n10115 ^ n10113 ;
  assign n10121 = n10119 & n10120 ;
  assign n10123 = n10121 ^ n10117 ;
  assign n10128 = n10125 ^ n10123 ;
  assign n10116 = n10111 ^ n10110 ;
  assign n10129 = n10128 ^ n10116 ;
  assign n10208 = n10161 ^ n10129 ;
  assign n10032 = n10027 ^ n10025 ;
  assign n10033 = n10028 ^ n10026 ;
  assign n10034 = n10032 & n10033 ;
  assign n10036 = n10034 ^ n10030 ;
  assign n10041 = n10038 ^ n10036 ;
  assign n10029 = n10024 ^ n10023 ;
  assign n10042 = n10041 ^ n10029 ;
  assign n10000 = n9995 ^ n9993 ;
  assign n10001 = n9996 ^ n9994 ;
  assign n10002 = n10000 & n10001 ;
  assign n10004 = n10002 ^ n9998 ;
  assign n10009 = n10006 ^ n10004 ;
  assign n9997 = n9992 ^ n9991 ;
  assign n10010 = n10009 ^ n9997 ;
  assign n10089 = n10042 ^ n10010 ;
  assign n10362 = n10208 ^ n10089 ;
  assign n11241 = n10766 ^ n10362 ;
  assign n9248 = n9243 ^ n9241 ;
  assign n9249 = n9244 ^ n9242 ;
  assign n9250 = n9248 & n9249 ;
  assign n9252 = n9250 ^ n9246 ;
  assign n9257 = n9254 ^ n9252 ;
  assign n9245 = n9240 ^ n9239 ;
  assign n9258 = n9257 ^ n9245 ;
  assign n9216 = n9211 ^ n9209 ;
  assign n9217 = n9212 ^ n9210 ;
  assign n9218 = n9216 & n9217 ;
  assign n9220 = n9218 ^ n9214 ;
  assign n9225 = n9222 ^ n9220 ;
  assign n9213 = n9208 ^ n9207 ;
  assign n9226 = n9225 ^ n9213 ;
  assign n9305 = n9258 ^ n9226 ;
  assign n9129 = n9124 ^ n9122 ;
  assign n9130 = n9125 ^ n9123 ;
  assign n9131 = n9129 & n9130 ;
  assign n9133 = n9131 ^ n9127 ;
  assign n9138 = n9135 ^ n9133 ;
  assign n9126 = n9121 ^ n9120 ;
  assign n9139 = n9138 ^ n9126 ;
  assign n9097 = n9092 ^ n9090 ;
  assign n9098 = n9093 ^ n9091 ;
  assign n9099 = n9097 & n9098 ;
  assign n9101 = n9099 ^ n9095 ;
  assign n9106 = n9103 ^ n9101 ;
  assign n9094 = n9089 ^ n9088 ;
  assign n9107 = n9106 ^ n9094 ;
  assign n9186 = n9139 ^ n9107 ;
  assign n9459 = n9305 ^ n9186 ;
  assign n8844 = n8839 ^ n8837 ;
  assign n8845 = n8840 ^ n8838 ;
  assign n8846 = n8844 & n8845 ;
  assign n8848 = n8846 ^ n8842 ;
  assign n8853 = n8850 ^ n8848 ;
  assign n8841 = n8836 ^ n8835 ;
  assign n8854 = n8853 ^ n8841 ;
  assign n8812 = n8807 ^ n8805 ;
  assign n8813 = n8808 ^ n8806 ;
  assign n8814 = n8812 & n8813 ;
  assign n8816 = n8814 ^ n8810 ;
  assign n8821 = n8818 ^ n8816 ;
  assign n8809 = n8804 ^ n8803 ;
  assign n8822 = n8821 ^ n8809 ;
  assign n8901 = n8854 ^ n8822 ;
  assign n8725 = n8720 ^ n8718 ;
  assign n8726 = n8721 ^ n8719 ;
  assign n8727 = n8725 & n8726 ;
  assign n8729 = n8727 ^ n8723 ;
  assign n8734 = n8731 ^ n8729 ;
  assign n8722 = n8717 ^ n8716 ;
  assign n8735 = n8734 ^ n8722 ;
  assign n8693 = n8688 ^ n8686 ;
  assign n8694 = n8689 ^ n8687 ;
  assign n8695 = n8693 & n8694 ;
  assign n8697 = n8695 ^ n8691 ;
  assign n8702 = n8699 ^ n8697 ;
  assign n8690 = n8685 ^ n8684 ;
  assign n8703 = n8702 ^ n8690 ;
  assign n8782 = n8735 ^ n8703 ;
  assign n9055 = n8901 ^ n8782 ;
  assign n9934 = n9459 ^ n9055 ;
  assign n12691 = n11241 ^ n9934 ;
  assign n12854 = n12787 ^ n12691 ;
  assign n12855 = n12854 ^ n8424 ;
  assign n10572 = n8607 ^ n8599 ;
  assign n10573 = n8608 ^ n8600 ;
  assign n10585 = n10572 & n10573 ;
  assign n10570 = n8605 ^ n8597 ;
  assign n10571 = n8606 ^ n8598 ;
  assign n10584 = n10570 & n10571 ;
  assign n10589 = n10585 ^ n10584 ;
  assign n10568 = n8603 ^ n8595 ;
  assign n10569 = n8604 ^ n8596 ;
  assign n10578 = n10568 & n10569 ;
  assign n10566 = n8601 ^ n8593 ;
  assign n10567 = n8602 ^ n8594 ;
  assign n10577 = n10566 & n10567 ;
  assign n10582 = n10578 ^ n10577 ;
  assign n10603 = n10589 ^ n10582 ;
  assign n10613 = n10609 ^ n10603 ;
  assign n10614 = n10613 ^ n10563 ;
  assign n10453 = n8591 ^ n8583 ;
  assign n10454 = n8592 ^ n8584 ;
  assign n10466 = n10453 & n10454 ;
  assign n10451 = n8589 ^ n8581 ;
  assign n10452 = n8590 ^ n8582 ;
  assign n10465 = n10451 & n10452 ;
  assign n10470 = n10466 ^ n10465 ;
  assign n10449 = n8587 ^ n8579 ;
  assign n10450 = n8588 ^ n8580 ;
  assign n10459 = n10449 & n10450 ;
  assign n10447 = n8585 ^ n8577 ;
  assign n10448 = n8586 ^ n8578 ;
  assign n10458 = n10447 & n10448 ;
  assign n10463 = n10459 ^ n10458 ;
  assign n10484 = n10470 ^ n10463 ;
  assign n10494 = n10490 ^ n10484 ;
  assign n10495 = n10494 ^ n10444 ;
  assign n10767 = n10614 ^ n10495 ;
  assign n10168 = n8575 ^ n8567 ;
  assign n10169 = n8576 ^ n8568 ;
  assign n10181 = n10168 & n10169 ;
  assign n10166 = n8573 ^ n8565 ;
  assign n10167 = n8574 ^ n8566 ;
  assign n10180 = n10166 & n10167 ;
  assign n10185 = n10181 ^ n10180 ;
  assign n10164 = n8571 ^ n8563 ;
  assign n10165 = n8572 ^ n8564 ;
  assign n10174 = n10164 & n10165 ;
  assign n10162 = n8569 ^ n8561 ;
  assign n10163 = n8570 ^ n8562 ;
  assign n10173 = n10162 & n10163 ;
  assign n10178 = n10174 ^ n10173 ;
  assign n10199 = n10185 ^ n10178 ;
  assign n10209 = n10205 ^ n10199 ;
  assign n10210 = n10209 ^ n10159 ;
  assign n10049 = n8559 ^ n8551 ;
  assign n10050 = n8560 ^ n8552 ;
  assign n10062 = n10049 & n10050 ;
  assign n10047 = n8557 ^ n8549 ;
  assign n10048 = n8558 ^ n8550 ;
  assign n10061 = n10047 & n10048 ;
  assign n10066 = n10062 ^ n10061 ;
  assign n10045 = n8555 ^ n8547 ;
  assign n10046 = n8556 ^ n8548 ;
  assign n10055 = n10045 & n10046 ;
  assign n10043 = n8553 ^ n8545 ;
  assign n10044 = n8554 ^ n8546 ;
  assign n10054 = n10043 & n10044 ;
  assign n10059 = n10055 ^ n10054 ;
  assign n10080 = n10066 ^ n10059 ;
  assign n10090 = n10086 ^ n10080 ;
  assign n10091 = n10090 ^ n10040 ;
  assign n10363 = n10210 ^ n10091 ;
  assign n11242 = n10767 ^ n10363 ;
  assign n9265 = n8543 ^ n8535 ;
  assign n9266 = n8544 ^ n8536 ;
  assign n9278 = n9265 & n9266 ;
  assign n9263 = n8541 ^ n8533 ;
  assign n9264 = n8542 ^ n8534 ;
  assign n9277 = n9263 & n9264 ;
  assign n9282 = n9278 ^ n9277 ;
  assign n9261 = n8539 ^ n8531 ;
  assign n9262 = n8540 ^ n8532 ;
  assign n9271 = n9261 & n9262 ;
  assign n9259 = n8537 ^ n8529 ;
  assign n9260 = n8538 ^ n8530 ;
  assign n9270 = n9259 & n9260 ;
  assign n9275 = n9271 ^ n9270 ;
  assign n9296 = n9282 ^ n9275 ;
  assign n9306 = n9302 ^ n9296 ;
  assign n9307 = n9306 ^ n9256 ;
  assign n9146 = n8527 ^ n8519 ;
  assign n9147 = n8528 ^ n8520 ;
  assign n9159 = n9146 & n9147 ;
  assign n9144 = n8525 ^ n8517 ;
  assign n9145 = n8526 ^ n8518 ;
  assign n9158 = n9144 & n9145 ;
  assign n9163 = n9159 ^ n9158 ;
  assign n9142 = n8523 ^ n8515 ;
  assign n9143 = n8524 ^ n8516 ;
  assign n9152 = n9142 & n9143 ;
  assign n9140 = n8521 ^ n8513 ;
  assign n9141 = n8522 ^ n8514 ;
  assign n9151 = n9140 & n9141 ;
  assign n9156 = n9152 ^ n9151 ;
  assign n9177 = n9163 ^ n9156 ;
  assign n9187 = n9183 ^ n9177 ;
  assign n9188 = n9187 ^ n9137 ;
  assign n9460 = n9307 ^ n9188 ;
  assign n8861 = n8511 ^ n8503 ;
  assign n8862 = n8512 ^ n8504 ;
  assign n8874 = n8861 & n8862 ;
  assign n8859 = n8509 ^ n8501 ;
  assign n8860 = n8510 ^ n8502 ;
  assign n8873 = n8859 & n8860 ;
  assign n8878 = n8874 ^ n8873 ;
  assign n8857 = n8507 ^ n8499 ;
  assign n8858 = n8508 ^ n8500 ;
  assign n8867 = n8857 & n8858 ;
  assign n8855 = n8505 ^ n8497 ;
  assign n8856 = n8506 ^ n8498 ;
  assign n8866 = n8855 & n8856 ;
  assign n8871 = n8867 ^ n8866 ;
  assign n8892 = n8878 ^ n8871 ;
  assign n8902 = n8898 ^ n8892 ;
  assign n8903 = n8902 ^ n8852 ;
  assign n8742 = n8495 ^ n8487 ;
  assign n8743 = n8496 ^ n8488 ;
  assign n8755 = n8742 & n8743 ;
  assign n8740 = n8493 ^ n8485 ;
  assign n8741 = n8494 ^ n8486 ;
  assign n8754 = n8740 & n8741 ;
  assign n8759 = n8755 ^ n8754 ;
  assign n8738 = n8491 ^ n8483 ;
  assign n8739 = n8492 ^ n8484 ;
  assign n8748 = n8738 & n8739 ;
  assign n8736 = n8489 ^ n8481 ;
  assign n8737 = n8490 ^ n8482 ;
  assign n8747 = n8736 & n8737 ;
  assign n8752 = n8748 ^ n8747 ;
  assign n8773 = n8759 ^ n8752 ;
  assign n8783 = n8779 ^ n8773 ;
  assign n8784 = n8783 ^ n8733 ;
  assign n9056 = n8903 ^ n8784 ;
  assign n9935 = n9460 ^ n9056 ;
  assign n12692 = n11242 ^ n9935 ;
  assign n12856 = n12788 ^ n12692 ;
  assign n12857 = n12856 ^ n8426 ;
  assign n10586 = n10572 ^ n10570 ;
  assign n10587 = n10573 ^ n10571 ;
  assign n10588 = n10586 & n10587 ;
  assign n10590 = n10588 ^ n10584 ;
  assign n10579 = n10568 ^ n10566 ;
  assign n10580 = n10569 ^ n10567 ;
  assign n10581 = n10579 & n10580 ;
  assign n10583 = n10581 ^ n10577 ;
  assign n10604 = n10590 ^ n10583 ;
  assign n10615 = n10610 ^ n10604 ;
  assign n10616 = n10615 ^ n10565 ;
  assign n10467 = n10453 ^ n10451 ;
  assign n10468 = n10454 ^ n10452 ;
  assign n10469 = n10467 & n10468 ;
  assign n10471 = n10469 ^ n10465 ;
  assign n10460 = n10449 ^ n10447 ;
  assign n10461 = n10450 ^ n10448 ;
  assign n10462 = n10460 & n10461 ;
  assign n10464 = n10462 ^ n10458 ;
  assign n10485 = n10471 ^ n10464 ;
  assign n10496 = n10491 ^ n10485 ;
  assign n10497 = n10496 ^ n10446 ;
  assign n10768 = n10616 ^ n10497 ;
  assign n10182 = n10168 ^ n10166 ;
  assign n10183 = n10169 ^ n10167 ;
  assign n10184 = n10182 & n10183 ;
  assign n10186 = n10184 ^ n10180 ;
  assign n10175 = n10164 ^ n10162 ;
  assign n10176 = n10165 ^ n10163 ;
  assign n10177 = n10175 & n10176 ;
  assign n10179 = n10177 ^ n10173 ;
  assign n10200 = n10186 ^ n10179 ;
  assign n10211 = n10206 ^ n10200 ;
  assign n10212 = n10211 ^ n10161 ;
  assign n10063 = n10049 ^ n10047 ;
  assign n10064 = n10050 ^ n10048 ;
  assign n10065 = n10063 & n10064 ;
  assign n10067 = n10065 ^ n10061 ;
  assign n10056 = n10045 ^ n10043 ;
  assign n10057 = n10046 ^ n10044 ;
  assign n10058 = n10056 & n10057 ;
  assign n10060 = n10058 ^ n10054 ;
  assign n10081 = n10067 ^ n10060 ;
  assign n10092 = n10087 ^ n10081 ;
  assign n10093 = n10092 ^ n10042 ;
  assign n10364 = n10212 ^ n10093 ;
  assign n11243 = n10768 ^ n10364 ;
  assign n9279 = n9265 ^ n9263 ;
  assign n9280 = n9266 ^ n9264 ;
  assign n9281 = n9279 & n9280 ;
  assign n9283 = n9281 ^ n9277 ;
  assign n9272 = n9261 ^ n9259 ;
  assign n9273 = n9262 ^ n9260 ;
  assign n9274 = n9272 & n9273 ;
  assign n9276 = n9274 ^ n9270 ;
  assign n9297 = n9283 ^ n9276 ;
  assign n9308 = n9303 ^ n9297 ;
  assign n9309 = n9308 ^ n9258 ;
  assign n9160 = n9146 ^ n9144 ;
  assign n9161 = n9147 ^ n9145 ;
  assign n9162 = n9160 & n9161 ;
  assign n9164 = n9162 ^ n9158 ;
  assign n9153 = n9142 ^ n9140 ;
  assign n9154 = n9143 ^ n9141 ;
  assign n9155 = n9153 & n9154 ;
  assign n9157 = n9155 ^ n9151 ;
  assign n9178 = n9164 ^ n9157 ;
  assign n9189 = n9184 ^ n9178 ;
  assign n9190 = n9189 ^ n9139 ;
  assign n9461 = n9309 ^ n9190 ;
  assign n8875 = n8861 ^ n8859 ;
  assign n8876 = n8862 ^ n8860 ;
  assign n8877 = n8875 & n8876 ;
  assign n8879 = n8877 ^ n8873 ;
  assign n8868 = n8857 ^ n8855 ;
  assign n8869 = n8858 ^ n8856 ;
  assign n8870 = n8868 & n8869 ;
  assign n8872 = n8870 ^ n8866 ;
  assign n8893 = n8879 ^ n8872 ;
  assign n8904 = n8899 ^ n8893 ;
  assign n8905 = n8904 ^ n8854 ;
  assign n8756 = n8742 ^ n8740 ;
  assign n8757 = n8743 ^ n8741 ;
  assign n8758 = n8756 & n8757 ;
  assign n8760 = n8758 ^ n8754 ;
  assign n8749 = n8738 ^ n8736 ;
  assign n8750 = n8739 ^ n8737 ;
  assign n8751 = n8749 & n8750 ;
  assign n8753 = n8751 ^ n8747 ;
  assign n8774 = n8760 ^ n8753 ;
  assign n8785 = n8780 ^ n8774 ;
  assign n8786 = n8785 ^ n8735 ;
  assign n9057 = n8905 ^ n8786 ;
  assign n9936 = n9461 ^ n9057 ;
  assign n12693 = n11243 ^ n9936 ;
  assign n12858 = n12789 ^ n12693 ;
  assign n12859 = n12858 ^ n8428 ;
  assign n10593 = n10572 ^ n10568 ;
  assign n10594 = n10573 ^ n10569 ;
  assign n10597 = n10593 & n10594 ;
  assign n10591 = n10570 ^ n10566 ;
  assign n10592 = n10571 ^ n10567 ;
  assign n10596 = n10591 & n10592 ;
  assign n10601 = n10597 ^ n10596 ;
  assign n10605 = n10603 ^ n10601 ;
  assign n10606 = n10605 ^ n10590 ;
  assign n10617 = n10611 ^ n10606 ;
  assign n10575 = n10565 ^ n10560 ;
  assign n10618 = n10617 ^ n10575 ;
  assign n10474 = n10453 ^ n10449 ;
  assign n10475 = n10454 ^ n10450 ;
  assign n10478 = n10474 & n10475 ;
  assign n10472 = n10451 ^ n10447 ;
  assign n10473 = n10452 ^ n10448 ;
  assign n10477 = n10472 & n10473 ;
  assign n10482 = n10478 ^ n10477 ;
  assign n10486 = n10484 ^ n10482 ;
  assign n10487 = n10486 ^ n10471 ;
  assign n10498 = n10492 ^ n10487 ;
  assign n10456 = n10446 ^ n10441 ;
  assign n10499 = n10498 ^ n10456 ;
  assign n10769 = n10618 ^ n10499 ;
  assign n10189 = n10168 ^ n10164 ;
  assign n10190 = n10169 ^ n10165 ;
  assign n10193 = n10189 & n10190 ;
  assign n10187 = n10166 ^ n10162 ;
  assign n10188 = n10167 ^ n10163 ;
  assign n10192 = n10187 & n10188 ;
  assign n10197 = n10193 ^ n10192 ;
  assign n10201 = n10199 ^ n10197 ;
  assign n10202 = n10201 ^ n10186 ;
  assign n10213 = n10207 ^ n10202 ;
  assign n10171 = n10161 ^ n10156 ;
  assign n10214 = n10213 ^ n10171 ;
  assign n10070 = n10049 ^ n10045 ;
  assign n10071 = n10050 ^ n10046 ;
  assign n10074 = n10070 & n10071 ;
  assign n10068 = n10047 ^ n10043 ;
  assign n10069 = n10048 ^ n10044 ;
  assign n10073 = n10068 & n10069 ;
  assign n10078 = n10074 ^ n10073 ;
  assign n10082 = n10080 ^ n10078 ;
  assign n10083 = n10082 ^ n10067 ;
  assign n10094 = n10088 ^ n10083 ;
  assign n10052 = n10042 ^ n10037 ;
  assign n10095 = n10094 ^ n10052 ;
  assign n10365 = n10214 ^ n10095 ;
  assign n11244 = n10769 ^ n10365 ;
  assign n9286 = n9265 ^ n9261 ;
  assign n9287 = n9266 ^ n9262 ;
  assign n9290 = n9286 & n9287 ;
  assign n9284 = n9263 ^ n9259 ;
  assign n9285 = n9264 ^ n9260 ;
  assign n9289 = n9284 & n9285 ;
  assign n9294 = n9290 ^ n9289 ;
  assign n9298 = n9296 ^ n9294 ;
  assign n9299 = n9298 ^ n9283 ;
  assign n9310 = n9304 ^ n9299 ;
  assign n9268 = n9258 ^ n9253 ;
  assign n9311 = n9310 ^ n9268 ;
  assign n9167 = n9146 ^ n9142 ;
  assign n9168 = n9147 ^ n9143 ;
  assign n9171 = n9167 & n9168 ;
  assign n9165 = n9144 ^ n9140 ;
  assign n9166 = n9145 ^ n9141 ;
  assign n9170 = n9165 & n9166 ;
  assign n9175 = n9171 ^ n9170 ;
  assign n9179 = n9177 ^ n9175 ;
  assign n9180 = n9179 ^ n9164 ;
  assign n9191 = n9185 ^ n9180 ;
  assign n9149 = n9139 ^ n9134 ;
  assign n9192 = n9191 ^ n9149 ;
  assign n9462 = n9311 ^ n9192 ;
  assign n8882 = n8861 ^ n8857 ;
  assign n8883 = n8862 ^ n8858 ;
  assign n8886 = n8882 & n8883 ;
  assign n8880 = n8859 ^ n8855 ;
  assign n8881 = n8860 ^ n8856 ;
  assign n8885 = n8880 & n8881 ;
  assign n8890 = n8886 ^ n8885 ;
  assign n8894 = n8892 ^ n8890 ;
  assign n8895 = n8894 ^ n8879 ;
  assign n8906 = n8900 ^ n8895 ;
  assign n8864 = n8854 ^ n8849 ;
  assign n8907 = n8906 ^ n8864 ;
  assign n8763 = n8742 ^ n8738 ;
  assign n8764 = n8743 ^ n8739 ;
  assign n8767 = n8763 & n8764 ;
  assign n8761 = n8740 ^ n8736 ;
  assign n8762 = n8741 ^ n8737 ;
  assign n8766 = n8761 & n8762 ;
  assign n8771 = n8767 ^ n8766 ;
  assign n8775 = n8773 ^ n8771 ;
  assign n8776 = n8775 ^ n8760 ;
  assign n8787 = n8781 ^ n8776 ;
  assign n8745 = n8735 ^ n8730 ;
  assign n8788 = n8787 ^ n8745 ;
  assign n9058 = n8907 ^ n8788 ;
  assign n9937 = n9462 ^ n9058 ;
  assign n12694 = n11244 ^ n9937 ;
  assign n12860 = n12790 ^ n12694 ;
  assign n12861 = n12860 ^ n8430 ;
  assign n10598 = n10593 ^ n10591 ;
  assign n10599 = n10594 ^ n10592 ;
  assign n10600 = n10598 & n10599 ;
  assign n10602 = n10600 ^ n10596 ;
  assign n10607 = n10604 ^ n10602 ;
  assign n10595 = n10590 ^ n10589 ;
  assign n10608 = n10607 ^ n10595 ;
  assign n10619 = n10612 ^ n10608 ;
  assign n10574 = n10565 ^ n10563 ;
  assign n10576 = n10574 ^ n10561 ;
  assign n10620 = n10619 ^ n10576 ;
  assign n10479 = n10474 ^ n10472 ;
  assign n10480 = n10475 ^ n10473 ;
  assign n10481 = n10479 & n10480 ;
  assign n10483 = n10481 ^ n10477 ;
  assign n10488 = n10485 ^ n10483 ;
  assign n10476 = n10471 ^ n10470 ;
  assign n10489 = n10488 ^ n10476 ;
  assign n10500 = n10493 ^ n10489 ;
  assign n10455 = n10446 ^ n10444 ;
  assign n10457 = n10455 ^ n10442 ;
  assign n10501 = n10500 ^ n10457 ;
  assign n10770 = n10620 ^ n10501 ;
  assign n10194 = n10189 ^ n10187 ;
  assign n10195 = n10190 ^ n10188 ;
  assign n10196 = n10194 & n10195 ;
  assign n10198 = n10196 ^ n10192 ;
  assign n10203 = n10200 ^ n10198 ;
  assign n10191 = n10186 ^ n10185 ;
  assign n10204 = n10203 ^ n10191 ;
  assign n10215 = n10208 ^ n10204 ;
  assign n10170 = n10161 ^ n10159 ;
  assign n10172 = n10170 ^ n10157 ;
  assign n10216 = n10215 ^ n10172 ;
  assign n10075 = n10070 ^ n10068 ;
  assign n10076 = n10071 ^ n10069 ;
  assign n10077 = n10075 & n10076 ;
  assign n10079 = n10077 ^ n10073 ;
  assign n10084 = n10081 ^ n10079 ;
  assign n10072 = n10067 ^ n10066 ;
  assign n10085 = n10084 ^ n10072 ;
  assign n10096 = n10089 ^ n10085 ;
  assign n10051 = n10042 ^ n10040 ;
  assign n10053 = n10051 ^ n10038 ;
  assign n10097 = n10096 ^ n10053 ;
  assign n10366 = n10216 ^ n10097 ;
  assign n11245 = n10770 ^ n10366 ;
  assign n9291 = n9286 ^ n9284 ;
  assign n9292 = n9287 ^ n9285 ;
  assign n9293 = n9291 & n9292 ;
  assign n9295 = n9293 ^ n9289 ;
  assign n9300 = n9297 ^ n9295 ;
  assign n9288 = n9283 ^ n9282 ;
  assign n9301 = n9300 ^ n9288 ;
  assign n9312 = n9305 ^ n9301 ;
  assign n9267 = n9258 ^ n9256 ;
  assign n9269 = n9267 ^ n9254 ;
  assign n9313 = n9312 ^ n9269 ;
  assign n9172 = n9167 ^ n9165 ;
  assign n9173 = n9168 ^ n9166 ;
  assign n9174 = n9172 & n9173 ;
  assign n9176 = n9174 ^ n9170 ;
  assign n9181 = n9178 ^ n9176 ;
  assign n9169 = n9164 ^ n9163 ;
  assign n9182 = n9181 ^ n9169 ;
  assign n9193 = n9186 ^ n9182 ;
  assign n9148 = n9139 ^ n9137 ;
  assign n9150 = n9148 ^ n9135 ;
  assign n9194 = n9193 ^ n9150 ;
  assign n9463 = n9313 ^ n9194 ;
  assign n8887 = n8882 ^ n8880 ;
  assign n8888 = n8883 ^ n8881 ;
  assign n8889 = n8887 & n8888 ;
  assign n8891 = n8889 ^ n8885 ;
  assign n8896 = n8893 ^ n8891 ;
  assign n8884 = n8879 ^ n8878 ;
  assign n8897 = n8896 ^ n8884 ;
  assign n8908 = n8901 ^ n8897 ;
  assign n8863 = n8854 ^ n8852 ;
  assign n8865 = n8863 ^ n8850 ;
  assign n8909 = n8908 ^ n8865 ;
  assign n8768 = n8763 ^ n8761 ;
  assign n8769 = n8764 ^ n8762 ;
  assign n8770 = n8768 & n8769 ;
  assign n8772 = n8770 ^ n8766 ;
  assign n8777 = n8774 ^ n8772 ;
  assign n8765 = n8760 ^ n8759 ;
  assign n8778 = n8777 ^ n8765 ;
  assign n8789 = n8782 ^ n8778 ;
  assign n8744 = n8735 ^ n8733 ;
  assign n8746 = n8744 ^ n8731 ;
  assign n8790 = n8789 ^ n8746 ;
  assign n9059 = n8909 ^ n8790 ;
  assign n9938 = n9463 ^ n9059 ;
  assign n12695 = n11245 ^ n9938 ;
  assign n12862 = n12791 ^ n12695 ;
  assign n12863 = n12862 ^ n8432 ;
  assign n10635 = n8607 ^ n8591 ;
  assign n10636 = n8608 ^ n8592 ;
  assign n10684 = n10635 & n10636 ;
  assign n10633 = n8605 ^ n8589 ;
  assign n10634 = n8606 ^ n8590 ;
  assign n10683 = n10633 & n10634 ;
  assign n10688 = n10684 ^ n10683 ;
  assign n10631 = n8603 ^ n8587 ;
  assign n10632 = n8604 ^ n8588 ;
  assign n10677 = n10631 & n10632 ;
  assign n10629 = n8601 ^ n8585 ;
  assign n10630 = n8602 ^ n8586 ;
  assign n10676 = n10629 & n10630 ;
  assign n10681 = n10677 ^ n10676 ;
  assign n10702 = n10688 ^ n10681 ;
  assign n10627 = n8599 ^ n8583 ;
  assign n10628 = n8600 ^ n8584 ;
  assign n10652 = n10627 & n10628 ;
  assign n10625 = n8597 ^ n8581 ;
  assign n10626 = n8598 ^ n8582 ;
  assign n10651 = n10625 & n10626 ;
  assign n10656 = n10652 ^ n10651 ;
  assign n10623 = n8595 ^ n8579 ;
  assign n10624 = n8596 ^ n8580 ;
  assign n10645 = n10623 & n10624 ;
  assign n10621 = n8593 ^ n8577 ;
  assign n10622 = n8594 ^ n8578 ;
  assign n10644 = n10621 & n10622 ;
  assign n10649 = n10645 ^ n10644 ;
  assign n10670 = n10656 ^ n10649 ;
  assign n10751 = n10702 ^ n10670 ;
  assign n10771 = n10763 ^ n10751 ;
  assign n10772 = n10771 ^ n10614 ;
  assign n10231 = n8575 ^ n8559 ;
  assign n10232 = n8576 ^ n8560 ;
  assign n10280 = n10231 & n10232 ;
  assign n10229 = n8573 ^ n8557 ;
  assign n10230 = n8574 ^ n8558 ;
  assign n10279 = n10229 & n10230 ;
  assign n10284 = n10280 ^ n10279 ;
  assign n10227 = n8571 ^ n8555 ;
  assign n10228 = n8572 ^ n8556 ;
  assign n10273 = n10227 & n10228 ;
  assign n10225 = n8569 ^ n8553 ;
  assign n10226 = n8570 ^ n8554 ;
  assign n10272 = n10225 & n10226 ;
  assign n10277 = n10273 ^ n10272 ;
  assign n10298 = n10284 ^ n10277 ;
  assign n10223 = n8567 ^ n8551 ;
  assign n10224 = n8568 ^ n8552 ;
  assign n10248 = n10223 & n10224 ;
  assign n10221 = n8565 ^ n8549 ;
  assign n10222 = n8566 ^ n8550 ;
  assign n10247 = n10221 & n10222 ;
  assign n10252 = n10248 ^ n10247 ;
  assign n10219 = n8563 ^ n8547 ;
  assign n10220 = n8564 ^ n8548 ;
  assign n10241 = n10219 & n10220 ;
  assign n10217 = n8561 ^ n8545 ;
  assign n10218 = n8562 ^ n8546 ;
  assign n10240 = n10217 & n10218 ;
  assign n10245 = n10241 ^ n10240 ;
  assign n10266 = n10252 ^ n10245 ;
  assign n10347 = n10298 ^ n10266 ;
  assign n10367 = n10359 ^ n10347 ;
  assign n10368 = n10367 ^ n10210 ;
  assign n11246 = n10772 ^ n10368 ;
  assign n9328 = n8543 ^ n8527 ;
  assign n9329 = n8544 ^ n8528 ;
  assign n9377 = n9328 & n9329 ;
  assign n9326 = n8541 ^ n8525 ;
  assign n9327 = n8542 ^ n8526 ;
  assign n9376 = n9326 & n9327 ;
  assign n9381 = n9377 ^ n9376 ;
  assign n9324 = n8539 ^ n8523 ;
  assign n9325 = n8540 ^ n8524 ;
  assign n9370 = n9324 & n9325 ;
  assign n9322 = n8537 ^ n8521 ;
  assign n9323 = n8538 ^ n8522 ;
  assign n9369 = n9322 & n9323 ;
  assign n9374 = n9370 ^ n9369 ;
  assign n9395 = n9381 ^ n9374 ;
  assign n9320 = n8535 ^ n8519 ;
  assign n9321 = n8536 ^ n8520 ;
  assign n9345 = n9320 & n9321 ;
  assign n9318 = n8533 ^ n8517 ;
  assign n9319 = n8534 ^ n8518 ;
  assign n9344 = n9318 & n9319 ;
  assign n9349 = n9345 ^ n9344 ;
  assign n9316 = n8531 ^ n8515 ;
  assign n9317 = n8532 ^ n8516 ;
  assign n9338 = n9316 & n9317 ;
  assign n9314 = n8529 ^ n8513 ;
  assign n9315 = n8530 ^ n8514 ;
  assign n9337 = n9314 & n9315 ;
  assign n9342 = n9338 ^ n9337 ;
  assign n9363 = n9349 ^ n9342 ;
  assign n9444 = n9395 ^ n9363 ;
  assign n9464 = n9456 ^ n9444 ;
  assign n9465 = n9464 ^ n9307 ;
  assign n8924 = n8511 ^ n8495 ;
  assign n8925 = n8512 ^ n8496 ;
  assign n8973 = n8924 & n8925 ;
  assign n8922 = n8509 ^ n8493 ;
  assign n8923 = n8510 ^ n8494 ;
  assign n8972 = n8922 & n8923 ;
  assign n8977 = n8973 ^ n8972 ;
  assign n8920 = n8507 ^ n8491 ;
  assign n8921 = n8508 ^ n8492 ;
  assign n8966 = n8920 & n8921 ;
  assign n8918 = n8505 ^ n8489 ;
  assign n8919 = n8506 ^ n8490 ;
  assign n8965 = n8918 & n8919 ;
  assign n8970 = n8966 ^ n8965 ;
  assign n8991 = n8977 ^ n8970 ;
  assign n8916 = n8503 ^ n8487 ;
  assign n8917 = n8504 ^ n8488 ;
  assign n8941 = n8916 & n8917 ;
  assign n8914 = n8501 ^ n8485 ;
  assign n8915 = n8502 ^ n8486 ;
  assign n8940 = n8914 & n8915 ;
  assign n8945 = n8941 ^ n8940 ;
  assign n8912 = n8499 ^ n8483 ;
  assign n8913 = n8500 ^ n8484 ;
  assign n8934 = n8912 & n8913 ;
  assign n8910 = n8497 ^ n8481 ;
  assign n8911 = n8498 ^ n8482 ;
  assign n8933 = n8910 & n8911 ;
  assign n8938 = n8934 ^ n8933 ;
  assign n8959 = n8945 ^ n8938 ;
  assign n9040 = n8991 ^ n8959 ;
  assign n9060 = n9052 ^ n9040 ;
  assign n9061 = n9060 ^ n8903 ;
  assign n9939 = n9465 ^ n9061 ;
  assign n12696 = n11246 ^ n9939 ;
  assign n12864 = n12792 ^ n12696 ;
  assign n12865 = n12864 ^ n8434 ;
  assign n10685 = n10635 ^ n10633 ;
  assign n10686 = n10636 ^ n10634 ;
  assign n10687 = n10685 & n10686 ;
  assign n10689 = n10687 ^ n10683 ;
  assign n10678 = n10631 ^ n10629 ;
  assign n10679 = n10632 ^ n10630 ;
  assign n10680 = n10678 & n10679 ;
  assign n10682 = n10680 ^ n10676 ;
  assign n10703 = n10689 ^ n10682 ;
  assign n10653 = n10627 ^ n10625 ;
  assign n10654 = n10628 ^ n10626 ;
  assign n10655 = n10653 & n10654 ;
  assign n10657 = n10655 ^ n10651 ;
  assign n10646 = n10623 ^ n10621 ;
  assign n10647 = n10624 ^ n10622 ;
  assign n10648 = n10646 & n10647 ;
  assign n10650 = n10648 ^ n10644 ;
  assign n10671 = n10657 ^ n10650 ;
  assign n10752 = n10703 ^ n10671 ;
  assign n10773 = n10764 ^ n10752 ;
  assign n10774 = n10773 ^ n10616 ;
  assign n10281 = n10231 ^ n10229 ;
  assign n10282 = n10232 ^ n10230 ;
  assign n10283 = n10281 & n10282 ;
  assign n10285 = n10283 ^ n10279 ;
  assign n10274 = n10227 ^ n10225 ;
  assign n10275 = n10228 ^ n10226 ;
  assign n10276 = n10274 & n10275 ;
  assign n10278 = n10276 ^ n10272 ;
  assign n10299 = n10285 ^ n10278 ;
  assign n10249 = n10223 ^ n10221 ;
  assign n10250 = n10224 ^ n10222 ;
  assign n10251 = n10249 & n10250 ;
  assign n10253 = n10251 ^ n10247 ;
  assign n10242 = n10219 ^ n10217 ;
  assign n10243 = n10220 ^ n10218 ;
  assign n10244 = n10242 & n10243 ;
  assign n10246 = n10244 ^ n10240 ;
  assign n10267 = n10253 ^ n10246 ;
  assign n10348 = n10299 ^ n10267 ;
  assign n10369 = n10360 ^ n10348 ;
  assign n10370 = n10369 ^ n10212 ;
  assign n11247 = n10774 ^ n10370 ;
  assign n9378 = n9328 ^ n9326 ;
  assign n9379 = n9329 ^ n9327 ;
  assign n9380 = n9378 & n9379 ;
  assign n9382 = n9380 ^ n9376 ;
  assign n9371 = n9324 ^ n9322 ;
  assign n9372 = n9325 ^ n9323 ;
  assign n9373 = n9371 & n9372 ;
  assign n9375 = n9373 ^ n9369 ;
  assign n9396 = n9382 ^ n9375 ;
  assign n9346 = n9320 ^ n9318 ;
  assign n9347 = n9321 ^ n9319 ;
  assign n9348 = n9346 & n9347 ;
  assign n9350 = n9348 ^ n9344 ;
  assign n9339 = n9316 ^ n9314 ;
  assign n9340 = n9317 ^ n9315 ;
  assign n9341 = n9339 & n9340 ;
  assign n9343 = n9341 ^ n9337 ;
  assign n9364 = n9350 ^ n9343 ;
  assign n9445 = n9396 ^ n9364 ;
  assign n9466 = n9457 ^ n9445 ;
  assign n9467 = n9466 ^ n9309 ;
  assign n8974 = n8924 ^ n8922 ;
  assign n8975 = n8925 ^ n8923 ;
  assign n8976 = n8974 & n8975 ;
  assign n8978 = n8976 ^ n8972 ;
  assign n8967 = n8920 ^ n8918 ;
  assign n8968 = n8921 ^ n8919 ;
  assign n8969 = n8967 & n8968 ;
  assign n8971 = n8969 ^ n8965 ;
  assign n8992 = n8978 ^ n8971 ;
  assign n8942 = n8916 ^ n8914 ;
  assign n8943 = n8917 ^ n8915 ;
  assign n8944 = n8942 & n8943 ;
  assign n8946 = n8944 ^ n8940 ;
  assign n8935 = n8912 ^ n8910 ;
  assign n8936 = n8913 ^ n8911 ;
  assign n8937 = n8935 & n8936 ;
  assign n8939 = n8937 ^ n8933 ;
  assign n8960 = n8946 ^ n8939 ;
  assign n9041 = n8992 ^ n8960 ;
  assign n9062 = n9053 ^ n9041 ;
  assign n9063 = n9062 ^ n8905 ;
  assign n9940 = n9467 ^ n9063 ;
  assign n12697 = n11247 ^ n9940 ;
  assign n12866 = n12793 ^ n12697 ;
  assign n12867 = n12866 ^ n8436 ;
  assign n10692 = n10635 ^ n10631 ;
  assign n10693 = n10636 ^ n10632 ;
  assign n10696 = n10692 & n10693 ;
  assign n10690 = n10633 ^ n10629 ;
  assign n10691 = n10634 ^ n10630 ;
  assign n10695 = n10690 & n10691 ;
  assign n10700 = n10696 ^ n10695 ;
  assign n10704 = n10702 ^ n10700 ;
  assign n10705 = n10704 ^ n10689 ;
  assign n10660 = n10627 ^ n10623 ;
  assign n10661 = n10628 ^ n10624 ;
  assign n10664 = n10660 & n10661 ;
  assign n10658 = n10625 ^ n10621 ;
  assign n10659 = n10626 ^ n10622 ;
  assign n10663 = n10658 & n10659 ;
  assign n10668 = n10664 ^ n10663 ;
  assign n10672 = n10670 ^ n10668 ;
  assign n10673 = n10672 ^ n10657 ;
  assign n10753 = n10705 ^ n10673 ;
  assign n10775 = n10765 ^ n10753 ;
  assign n10776 = n10775 ^ n10618 ;
  assign n10288 = n10231 ^ n10227 ;
  assign n10289 = n10232 ^ n10228 ;
  assign n10292 = n10288 & n10289 ;
  assign n10286 = n10229 ^ n10225 ;
  assign n10287 = n10230 ^ n10226 ;
  assign n10291 = n10286 & n10287 ;
  assign n10296 = n10292 ^ n10291 ;
  assign n10300 = n10298 ^ n10296 ;
  assign n10301 = n10300 ^ n10285 ;
  assign n10256 = n10223 ^ n10219 ;
  assign n10257 = n10224 ^ n10220 ;
  assign n10260 = n10256 & n10257 ;
  assign n10254 = n10221 ^ n10217 ;
  assign n10255 = n10222 ^ n10218 ;
  assign n10259 = n10254 & n10255 ;
  assign n10264 = n10260 ^ n10259 ;
  assign n10268 = n10266 ^ n10264 ;
  assign n10269 = n10268 ^ n10253 ;
  assign n10349 = n10301 ^ n10269 ;
  assign n10371 = n10361 ^ n10349 ;
  assign n10372 = n10371 ^ n10214 ;
  assign n11248 = n10776 ^ n10372 ;
  assign n9385 = n9328 ^ n9324 ;
  assign n9386 = n9329 ^ n9325 ;
  assign n9389 = n9385 & n9386 ;
  assign n9383 = n9326 ^ n9322 ;
  assign n9384 = n9327 ^ n9323 ;
  assign n9388 = n9383 & n9384 ;
  assign n9393 = n9389 ^ n9388 ;
  assign n9397 = n9395 ^ n9393 ;
  assign n9398 = n9397 ^ n9382 ;
  assign n9353 = n9320 ^ n9316 ;
  assign n9354 = n9321 ^ n9317 ;
  assign n9357 = n9353 & n9354 ;
  assign n9351 = n9318 ^ n9314 ;
  assign n9352 = n9319 ^ n9315 ;
  assign n9356 = n9351 & n9352 ;
  assign n9361 = n9357 ^ n9356 ;
  assign n9365 = n9363 ^ n9361 ;
  assign n9366 = n9365 ^ n9350 ;
  assign n9446 = n9398 ^ n9366 ;
  assign n9468 = n9458 ^ n9446 ;
  assign n9469 = n9468 ^ n9311 ;
  assign n8981 = n8924 ^ n8920 ;
  assign n8982 = n8925 ^ n8921 ;
  assign n8985 = n8981 & n8982 ;
  assign n8979 = n8922 ^ n8918 ;
  assign n8980 = n8923 ^ n8919 ;
  assign n8984 = n8979 & n8980 ;
  assign n8989 = n8985 ^ n8984 ;
  assign n8993 = n8991 ^ n8989 ;
  assign n8994 = n8993 ^ n8978 ;
  assign n8949 = n8916 ^ n8912 ;
  assign n8950 = n8917 ^ n8913 ;
  assign n8953 = n8949 & n8950 ;
  assign n8947 = n8914 ^ n8910 ;
  assign n8948 = n8915 ^ n8911 ;
  assign n8952 = n8947 & n8948 ;
  assign n8957 = n8953 ^ n8952 ;
  assign n8961 = n8959 ^ n8957 ;
  assign n8962 = n8961 ^ n8946 ;
  assign n9042 = n8994 ^ n8962 ;
  assign n9064 = n9054 ^ n9042 ;
  assign n9065 = n9064 ^ n8907 ;
  assign n9941 = n9469 ^ n9065 ;
  assign n12698 = n11248 ^ n9941 ;
  assign n12868 = n12794 ^ n12698 ;
  assign n12869 = n12868 ^ n8438 ;
  assign n10697 = n10692 ^ n10690 ;
  assign n10698 = n10693 ^ n10691 ;
  assign n10699 = n10697 & n10698 ;
  assign n10701 = n10699 ^ n10695 ;
  assign n10706 = n10703 ^ n10701 ;
  assign n10694 = n10689 ^ n10688 ;
  assign n10707 = n10706 ^ n10694 ;
  assign n10665 = n10660 ^ n10658 ;
  assign n10666 = n10661 ^ n10659 ;
  assign n10667 = n10665 & n10666 ;
  assign n10669 = n10667 ^ n10663 ;
  assign n10674 = n10671 ^ n10669 ;
  assign n10662 = n10657 ^ n10656 ;
  assign n10675 = n10674 ^ n10662 ;
  assign n10754 = n10707 ^ n10675 ;
  assign n10777 = n10766 ^ n10754 ;
  assign n10778 = n10777 ^ n10620 ;
  assign n10293 = n10288 ^ n10286 ;
  assign n10294 = n10289 ^ n10287 ;
  assign n10295 = n10293 & n10294 ;
  assign n10297 = n10295 ^ n10291 ;
  assign n10302 = n10299 ^ n10297 ;
  assign n10290 = n10285 ^ n10284 ;
  assign n10303 = n10302 ^ n10290 ;
  assign n10261 = n10256 ^ n10254 ;
  assign n10262 = n10257 ^ n10255 ;
  assign n10263 = n10261 & n10262 ;
  assign n10265 = n10263 ^ n10259 ;
  assign n10270 = n10267 ^ n10265 ;
  assign n10258 = n10253 ^ n10252 ;
  assign n10271 = n10270 ^ n10258 ;
  assign n10350 = n10303 ^ n10271 ;
  assign n10373 = n10362 ^ n10350 ;
  assign n10374 = n10373 ^ n10216 ;
  assign n11249 = n10778 ^ n10374 ;
  assign n9390 = n9385 ^ n9383 ;
  assign n9391 = n9386 ^ n9384 ;
  assign n9392 = n9390 & n9391 ;
  assign n9394 = n9392 ^ n9388 ;
  assign n9399 = n9396 ^ n9394 ;
  assign n9387 = n9382 ^ n9381 ;
  assign n9400 = n9399 ^ n9387 ;
  assign n9358 = n9353 ^ n9351 ;
  assign n9359 = n9354 ^ n9352 ;
  assign n9360 = n9358 & n9359 ;
  assign n9362 = n9360 ^ n9356 ;
  assign n9367 = n9364 ^ n9362 ;
  assign n9355 = n9350 ^ n9349 ;
  assign n9368 = n9367 ^ n9355 ;
  assign n9447 = n9400 ^ n9368 ;
  assign n9470 = n9459 ^ n9447 ;
  assign n9471 = n9470 ^ n9313 ;
  assign n8986 = n8981 ^ n8979 ;
  assign n8987 = n8982 ^ n8980 ;
  assign n8988 = n8986 & n8987 ;
  assign n8990 = n8988 ^ n8984 ;
  assign n8995 = n8992 ^ n8990 ;
  assign n8983 = n8978 ^ n8977 ;
  assign n8996 = n8995 ^ n8983 ;
  assign n8954 = n8949 ^ n8947 ;
  assign n8955 = n8950 ^ n8948 ;
  assign n8956 = n8954 & n8955 ;
  assign n8958 = n8956 ^ n8952 ;
  assign n8963 = n8960 ^ n8958 ;
  assign n8951 = n8946 ^ n8945 ;
  assign n8964 = n8963 ^ n8951 ;
  assign n9043 = n8996 ^ n8964 ;
  assign n9066 = n9055 ^ n9043 ;
  assign n9067 = n9066 ^ n8909 ;
  assign n9942 = n9471 ^ n9067 ;
  assign n12699 = n11249 ^ n9942 ;
  assign n12870 = n12795 ^ n12699 ;
  assign n12871 = n12870 ^ n8440 ;
  assign n10714 = n10635 ^ n10627 ;
  assign n10715 = n10636 ^ n10628 ;
  assign n10727 = n10714 & n10715 ;
  assign n10712 = n10633 ^ n10625 ;
  assign n10713 = n10634 ^ n10626 ;
  assign n10726 = n10712 & n10713 ;
  assign n10731 = n10727 ^ n10726 ;
  assign n10710 = n10631 ^ n10623 ;
  assign n10711 = n10632 ^ n10624 ;
  assign n10720 = n10710 & n10711 ;
  assign n10708 = n10629 ^ n10621 ;
  assign n10709 = n10630 ^ n10622 ;
  assign n10719 = n10708 & n10709 ;
  assign n10724 = n10720 ^ n10719 ;
  assign n10745 = n10731 ^ n10724 ;
  assign n10755 = n10751 ^ n10745 ;
  assign n10756 = n10755 ^ n10705 ;
  assign n10779 = n10767 ^ n10756 ;
  assign n10640 = n10618 ^ n10609 ;
  assign n10780 = n10779 ^ n10640 ;
  assign n10310 = n10231 ^ n10223 ;
  assign n10311 = n10232 ^ n10224 ;
  assign n10323 = n10310 & n10311 ;
  assign n10308 = n10229 ^ n10221 ;
  assign n10309 = n10230 ^ n10222 ;
  assign n10322 = n10308 & n10309 ;
  assign n10327 = n10323 ^ n10322 ;
  assign n10306 = n10227 ^ n10219 ;
  assign n10307 = n10228 ^ n10220 ;
  assign n10316 = n10306 & n10307 ;
  assign n10304 = n10225 ^ n10217 ;
  assign n10305 = n10226 ^ n10218 ;
  assign n10315 = n10304 & n10305 ;
  assign n10320 = n10316 ^ n10315 ;
  assign n10341 = n10327 ^ n10320 ;
  assign n10351 = n10347 ^ n10341 ;
  assign n10352 = n10351 ^ n10301 ;
  assign n10375 = n10363 ^ n10352 ;
  assign n10236 = n10214 ^ n10205 ;
  assign n10376 = n10375 ^ n10236 ;
  assign n11250 = n10780 ^ n10376 ;
  assign n9407 = n9328 ^ n9320 ;
  assign n9408 = n9329 ^ n9321 ;
  assign n9420 = n9407 & n9408 ;
  assign n9405 = n9326 ^ n9318 ;
  assign n9406 = n9327 ^ n9319 ;
  assign n9419 = n9405 & n9406 ;
  assign n9424 = n9420 ^ n9419 ;
  assign n9403 = n9324 ^ n9316 ;
  assign n9404 = n9325 ^ n9317 ;
  assign n9413 = n9403 & n9404 ;
  assign n9401 = n9322 ^ n9314 ;
  assign n9402 = n9323 ^ n9315 ;
  assign n9412 = n9401 & n9402 ;
  assign n9417 = n9413 ^ n9412 ;
  assign n9438 = n9424 ^ n9417 ;
  assign n9448 = n9444 ^ n9438 ;
  assign n9449 = n9448 ^ n9398 ;
  assign n9472 = n9460 ^ n9449 ;
  assign n9333 = n9311 ^ n9302 ;
  assign n9473 = n9472 ^ n9333 ;
  assign n9003 = n8924 ^ n8916 ;
  assign n9004 = n8925 ^ n8917 ;
  assign n9016 = n9003 & n9004 ;
  assign n9001 = n8922 ^ n8914 ;
  assign n9002 = n8923 ^ n8915 ;
  assign n9015 = n9001 & n9002 ;
  assign n9020 = n9016 ^ n9015 ;
  assign n8999 = n8920 ^ n8912 ;
  assign n9000 = n8921 ^ n8913 ;
  assign n9009 = n8999 & n9000 ;
  assign n8997 = n8918 ^ n8910 ;
  assign n8998 = n8919 ^ n8911 ;
  assign n9008 = n8997 & n8998 ;
  assign n9013 = n9009 ^ n9008 ;
  assign n9034 = n9020 ^ n9013 ;
  assign n9044 = n9040 ^ n9034 ;
  assign n9045 = n9044 ^ n8994 ;
  assign n9068 = n9056 ^ n9045 ;
  assign n8929 = n8907 ^ n8898 ;
  assign n9069 = n9068 ^ n8929 ;
  assign n9943 = n9473 ^ n9069 ;
  assign n12700 = n11250 ^ n9943 ;
  assign n12872 = n12796 ^ n12700 ;
  assign n12873 = n12872 ^ n8442 ;
  assign n10728 = n10714 ^ n10712 ;
  assign n10729 = n10715 ^ n10713 ;
  assign n10730 = n10728 & n10729 ;
  assign n10732 = n10730 ^ n10726 ;
  assign n10721 = n10710 ^ n10708 ;
  assign n10722 = n10711 ^ n10709 ;
  assign n10723 = n10721 & n10722 ;
  assign n10725 = n10723 ^ n10719 ;
  assign n10746 = n10732 ^ n10725 ;
  assign n10757 = n10752 ^ n10746 ;
  assign n10758 = n10757 ^ n10707 ;
  assign n10781 = n10768 ^ n10758 ;
  assign n10641 = n10620 ^ n10610 ;
  assign n10782 = n10781 ^ n10641 ;
  assign n10324 = n10310 ^ n10308 ;
  assign n10325 = n10311 ^ n10309 ;
  assign n10326 = n10324 & n10325 ;
  assign n10328 = n10326 ^ n10322 ;
  assign n10317 = n10306 ^ n10304 ;
  assign n10318 = n10307 ^ n10305 ;
  assign n10319 = n10317 & n10318 ;
  assign n10321 = n10319 ^ n10315 ;
  assign n10342 = n10328 ^ n10321 ;
  assign n10353 = n10348 ^ n10342 ;
  assign n10354 = n10353 ^ n10303 ;
  assign n10377 = n10364 ^ n10354 ;
  assign n10237 = n10216 ^ n10206 ;
  assign n10378 = n10377 ^ n10237 ;
  assign n11251 = n10782 ^ n10378 ;
  assign n9421 = n9407 ^ n9405 ;
  assign n9422 = n9408 ^ n9406 ;
  assign n9423 = n9421 & n9422 ;
  assign n9425 = n9423 ^ n9419 ;
  assign n9414 = n9403 ^ n9401 ;
  assign n9415 = n9404 ^ n9402 ;
  assign n9416 = n9414 & n9415 ;
  assign n9418 = n9416 ^ n9412 ;
  assign n9439 = n9425 ^ n9418 ;
  assign n9450 = n9445 ^ n9439 ;
  assign n9451 = n9450 ^ n9400 ;
  assign n9474 = n9461 ^ n9451 ;
  assign n9334 = n9313 ^ n9303 ;
  assign n9475 = n9474 ^ n9334 ;
  assign n9017 = n9003 ^ n9001 ;
  assign n9018 = n9004 ^ n9002 ;
  assign n9019 = n9017 & n9018 ;
  assign n9021 = n9019 ^ n9015 ;
  assign n9010 = n8999 ^ n8997 ;
  assign n9011 = n9000 ^ n8998 ;
  assign n9012 = n9010 & n9011 ;
  assign n9014 = n9012 ^ n9008 ;
  assign n9035 = n9021 ^ n9014 ;
  assign n9046 = n9041 ^ n9035 ;
  assign n9047 = n9046 ^ n8996 ;
  assign n9070 = n9057 ^ n9047 ;
  assign n8930 = n8909 ^ n8899 ;
  assign n9071 = n9070 ^ n8930 ;
  assign n9944 = n9475 ^ n9071 ;
  assign n12701 = n11251 ^ n9944 ;
  assign n12874 = n12797 ^ n12701 ;
  assign n12875 = n12874 ^ n8444 ;
  assign n10735 = n10714 ^ n10710 ;
  assign n10736 = n10715 ^ n10711 ;
  assign n10739 = n10735 & n10736 ;
  assign n10733 = n10712 ^ n10708 ;
  assign n10734 = n10713 ^ n10709 ;
  assign n10738 = n10733 & n10734 ;
  assign n10743 = n10739 ^ n10738 ;
  assign n10747 = n10745 ^ n10743 ;
  assign n10748 = n10747 ^ n10732 ;
  assign n10759 = n10753 ^ n10748 ;
  assign n10717 = n10707 ^ n10702 ;
  assign n10760 = n10759 ^ n10717 ;
  assign n10783 = n10769 ^ n10760 ;
  assign n10638 = n10620 ^ n10614 ;
  assign n10642 = n10638 ^ n10611 ;
  assign n10784 = n10783 ^ n10642 ;
  assign n10331 = n10310 ^ n10306 ;
  assign n10332 = n10311 ^ n10307 ;
  assign n10335 = n10331 & n10332 ;
  assign n10329 = n10308 ^ n10304 ;
  assign n10330 = n10309 ^ n10305 ;
  assign n10334 = n10329 & n10330 ;
  assign n10339 = n10335 ^ n10334 ;
  assign n10343 = n10341 ^ n10339 ;
  assign n10344 = n10343 ^ n10328 ;
  assign n10355 = n10349 ^ n10344 ;
  assign n10313 = n10303 ^ n10298 ;
  assign n10356 = n10355 ^ n10313 ;
  assign n10379 = n10365 ^ n10356 ;
  assign n10234 = n10216 ^ n10210 ;
  assign n10238 = n10234 ^ n10207 ;
  assign n10380 = n10379 ^ n10238 ;
  assign n11252 = n10784 ^ n10380 ;
  assign n9428 = n9407 ^ n9403 ;
  assign n9429 = n9408 ^ n9404 ;
  assign n9432 = n9428 & n9429 ;
  assign n9426 = n9405 ^ n9401 ;
  assign n9427 = n9406 ^ n9402 ;
  assign n9431 = n9426 & n9427 ;
  assign n9436 = n9432 ^ n9431 ;
  assign n9440 = n9438 ^ n9436 ;
  assign n9441 = n9440 ^ n9425 ;
  assign n9452 = n9446 ^ n9441 ;
  assign n9410 = n9400 ^ n9395 ;
  assign n9453 = n9452 ^ n9410 ;
  assign n9476 = n9462 ^ n9453 ;
  assign n9331 = n9313 ^ n9307 ;
  assign n9335 = n9331 ^ n9304 ;
  assign n9477 = n9476 ^ n9335 ;
  assign n9024 = n9003 ^ n8999 ;
  assign n9025 = n9004 ^ n9000 ;
  assign n9028 = n9024 & n9025 ;
  assign n9022 = n9001 ^ n8997 ;
  assign n9023 = n9002 ^ n8998 ;
  assign n9027 = n9022 & n9023 ;
  assign n9032 = n9028 ^ n9027 ;
  assign n9036 = n9034 ^ n9032 ;
  assign n9037 = n9036 ^ n9021 ;
  assign n9048 = n9042 ^ n9037 ;
  assign n9006 = n8996 ^ n8991 ;
  assign n9049 = n9048 ^ n9006 ;
  assign n9072 = n9058 ^ n9049 ;
  assign n8927 = n8909 ^ n8903 ;
  assign n8931 = n8927 ^ n8900 ;
  assign n9073 = n9072 ^ n8931 ;
  assign n9945 = n9477 ^ n9073 ;
  assign n12702 = n11252 ^ n9945 ;
  assign n12876 = n12798 ^ n12702 ;
  assign n12877 = n12876 ^ n8446 ;
  assign n10740 = n10735 ^ n10733 ;
  assign n10741 = n10736 ^ n10734 ;
  assign n10742 = n10740 & n10741 ;
  assign n10744 = n10742 ^ n10738 ;
  assign n10749 = n10746 ^ n10744 ;
  assign n10737 = n10732 ^ n10731 ;
  assign n10750 = n10749 ^ n10737 ;
  assign n10761 = n10754 ^ n10750 ;
  assign n10716 = n10707 ^ n10705 ;
  assign n10718 = n10716 ^ n10703 ;
  assign n10762 = n10761 ^ n10718 ;
  assign n10785 = n10770 ^ n10762 ;
  assign n10637 = n10620 ^ n10618 ;
  assign n10639 = n10637 ^ n10616 ;
  assign n10643 = n10639 ^ n10612 ;
  assign n10786 = n10785 ^ n10643 ;
  assign n10336 = n10331 ^ n10329 ;
  assign n10337 = n10332 ^ n10330 ;
  assign n10338 = n10336 & n10337 ;
  assign n10340 = n10338 ^ n10334 ;
  assign n10345 = n10342 ^ n10340 ;
  assign n10333 = n10328 ^ n10327 ;
  assign n10346 = n10345 ^ n10333 ;
  assign n10357 = n10350 ^ n10346 ;
  assign n10312 = n10303 ^ n10301 ;
  assign n10314 = n10312 ^ n10299 ;
  assign n10358 = n10357 ^ n10314 ;
  assign n10381 = n10366 ^ n10358 ;
  assign n10233 = n10216 ^ n10214 ;
  assign n10235 = n10233 ^ n10212 ;
  assign n10239 = n10235 ^ n10208 ;
  assign n10382 = n10381 ^ n10239 ;
  assign n11253 = n10786 ^ n10382 ;
  assign n9433 = n9428 ^ n9426 ;
  assign n9434 = n9429 ^ n9427 ;
  assign n9435 = n9433 & n9434 ;
  assign n9437 = n9435 ^ n9431 ;
  assign n9442 = n9439 ^ n9437 ;
  assign n9430 = n9425 ^ n9424 ;
  assign n9443 = n9442 ^ n9430 ;
  assign n9454 = n9447 ^ n9443 ;
  assign n9409 = n9400 ^ n9398 ;
  assign n9411 = n9409 ^ n9396 ;
  assign n9455 = n9454 ^ n9411 ;
  assign n9478 = n9463 ^ n9455 ;
  assign n9330 = n9313 ^ n9311 ;
  assign n9332 = n9330 ^ n9309 ;
  assign n9336 = n9332 ^ n9305 ;
  assign n9479 = n9478 ^ n9336 ;
  assign n9029 = n9024 ^ n9022 ;
  assign n9030 = n9025 ^ n9023 ;
  assign n9031 = n9029 & n9030 ;
  assign n9033 = n9031 ^ n9027 ;
  assign n9038 = n9035 ^ n9033 ;
  assign n9026 = n9021 ^ n9020 ;
  assign n9039 = n9038 ^ n9026 ;
  assign n9050 = n9043 ^ n9039 ;
  assign n9005 = n8996 ^ n8994 ;
  assign n9007 = n9005 ^ n8992 ;
  assign n9051 = n9050 ^ n9007 ;
  assign n9074 = n9059 ^ n9051 ;
  assign n8926 = n8909 ^ n8907 ;
  assign n8928 = n8926 ^ n8905 ;
  assign n8932 = n8928 ^ n8901 ;
  assign n9075 = n9074 ^ n8932 ;
  assign n9946 = n9479 ^ n9075 ;
  assign n12703 = n11253 ^ n9946 ;
  assign n12878 = n12799 ^ n12703 ;
  assign n12879 = n12878 ^ n8448 ;
  assign n10817 = n8607 ^ n8575 ;
  assign n10818 = n8608 ^ n8576 ;
  assign n10993 = n10817 & n10818 ;
  assign n10815 = n8605 ^ n8573 ;
  assign n10816 = n8606 ^ n8574 ;
  assign n10992 = n10815 & n10816 ;
  assign n10997 = n10993 ^ n10992 ;
  assign n10813 = n8603 ^ n8571 ;
  assign n10814 = n8604 ^ n8572 ;
  assign n10986 = n10813 & n10814 ;
  assign n10811 = n8601 ^ n8569 ;
  assign n10812 = n8602 ^ n8570 ;
  assign n10985 = n10811 & n10812 ;
  assign n10990 = n10986 ^ n10985 ;
  assign n11011 = n10997 ^ n10990 ;
  assign n10809 = n8599 ^ n8567 ;
  assign n10810 = n8600 ^ n8568 ;
  assign n10961 = n10809 & n10810 ;
  assign n10807 = n8597 ^ n8565 ;
  assign n10808 = n8598 ^ n8566 ;
  assign n10960 = n10807 & n10808 ;
  assign n10965 = n10961 ^ n10960 ;
  assign n10805 = n8595 ^ n8563 ;
  assign n10806 = n8596 ^ n8564 ;
  assign n10954 = n10805 & n10806 ;
  assign n10803 = n8593 ^ n8561 ;
  assign n10804 = n8594 ^ n8562 ;
  assign n10953 = n10803 & n10804 ;
  assign n10958 = n10954 ^ n10953 ;
  assign n10979 = n10965 ^ n10958 ;
  assign n11060 = n11011 ^ n10979 ;
  assign n10801 = n8591 ^ n8559 ;
  assign n10802 = n8592 ^ n8560 ;
  assign n10874 = n10801 & n10802 ;
  assign n10799 = n8589 ^ n8557 ;
  assign n10800 = n8590 ^ n8558 ;
  assign n10873 = n10799 & n10800 ;
  assign n10878 = n10874 ^ n10873 ;
  assign n10797 = n8587 ^ n8555 ;
  assign n10798 = n8588 ^ n8556 ;
  assign n10867 = n10797 & n10798 ;
  assign n10795 = n8585 ^ n8553 ;
  assign n10796 = n8586 ^ n8554 ;
  assign n10866 = n10795 & n10796 ;
  assign n10871 = n10867 ^ n10866 ;
  assign n10892 = n10878 ^ n10871 ;
  assign n10793 = n8583 ^ n8551 ;
  assign n10794 = n8584 ^ n8552 ;
  assign n10842 = n10793 & n10794 ;
  assign n10791 = n8581 ^ n8549 ;
  assign n10792 = n8582 ^ n8550 ;
  assign n10841 = n10791 & n10792 ;
  assign n10846 = n10842 ^ n10841 ;
  assign n10789 = n8579 ^ n8547 ;
  assign n10790 = n8580 ^ n8548 ;
  assign n10835 = n10789 & n10790 ;
  assign n10787 = n8577 ^ n8545 ;
  assign n10788 = n8578 ^ n8546 ;
  assign n10834 = n10787 & n10788 ;
  assign n10839 = n10835 ^ n10834 ;
  assign n10860 = n10846 ^ n10839 ;
  assign n10941 = n10892 ^ n10860 ;
  assign n11214 = n11060 ^ n10941 ;
  assign n11254 = n11238 ^ n11214 ;
  assign n11255 = n11254 ^ n10772 ;
  assign n9510 = n8543 ^ n8511 ;
  assign n9511 = n8544 ^ n8512 ;
  assign n9686 = n9510 & n9511 ;
  assign n9508 = n8541 ^ n8509 ;
  assign n9509 = n8542 ^ n8510 ;
  assign n9685 = n9508 & n9509 ;
  assign n9690 = n9686 ^ n9685 ;
  assign n9506 = n8539 ^ n8507 ;
  assign n9507 = n8540 ^ n8508 ;
  assign n9679 = n9506 & n9507 ;
  assign n9504 = n8537 ^ n8505 ;
  assign n9505 = n8538 ^ n8506 ;
  assign n9678 = n9504 & n9505 ;
  assign n9683 = n9679 ^ n9678 ;
  assign n9704 = n9690 ^ n9683 ;
  assign n9502 = n8535 ^ n8503 ;
  assign n9503 = n8536 ^ n8504 ;
  assign n9654 = n9502 & n9503 ;
  assign n9500 = n8533 ^ n8501 ;
  assign n9501 = n8534 ^ n8502 ;
  assign n9653 = n9500 & n9501 ;
  assign n9658 = n9654 ^ n9653 ;
  assign n9498 = n8531 ^ n8499 ;
  assign n9499 = n8532 ^ n8500 ;
  assign n9647 = n9498 & n9499 ;
  assign n9496 = n8529 ^ n8497 ;
  assign n9497 = n8530 ^ n8498 ;
  assign n9646 = n9496 & n9497 ;
  assign n9651 = n9647 ^ n9646 ;
  assign n9672 = n9658 ^ n9651 ;
  assign n9753 = n9704 ^ n9672 ;
  assign n9494 = n8527 ^ n8495 ;
  assign n9495 = n8528 ^ n8496 ;
  assign n9567 = n9494 & n9495 ;
  assign n9492 = n8525 ^ n8493 ;
  assign n9493 = n8526 ^ n8494 ;
  assign n9566 = n9492 & n9493 ;
  assign n9571 = n9567 ^ n9566 ;
  assign n9490 = n8523 ^ n8491 ;
  assign n9491 = n8524 ^ n8492 ;
  assign n9560 = n9490 & n9491 ;
  assign n9488 = n8521 ^ n8489 ;
  assign n9489 = n8522 ^ n8490 ;
  assign n9559 = n9488 & n9489 ;
  assign n9564 = n9560 ^ n9559 ;
  assign n9585 = n9571 ^ n9564 ;
  assign n9486 = n8519 ^ n8487 ;
  assign n9487 = n8520 ^ n8488 ;
  assign n9535 = n9486 & n9487 ;
  assign n9484 = n8517 ^ n8485 ;
  assign n9485 = n8518 ^ n8486 ;
  assign n9534 = n9484 & n9485 ;
  assign n9539 = n9535 ^ n9534 ;
  assign n9482 = n8515 ^ n8483 ;
  assign n9483 = n8516 ^ n8484 ;
  assign n9528 = n9482 & n9483 ;
  assign n9480 = n8513 ^ n8481 ;
  assign n9481 = n8514 ^ n8482 ;
  assign n9527 = n9480 & n9481 ;
  assign n9532 = n9528 ^ n9527 ;
  assign n9553 = n9539 ^ n9532 ;
  assign n9634 = n9585 ^ n9553 ;
  assign n9907 = n9753 ^ n9634 ;
  assign n9947 = n9931 ^ n9907 ;
  assign n9948 = n9947 ^ n9465 ;
  assign n12704 = n11255 ^ n9948 ;
  assign n12880 = n12800 ^ n12704 ;
  assign n12881 = n12880 ^ n8450 ;
  assign n10994 = n10817 ^ n10815 ;
  assign n10995 = n10818 ^ n10816 ;
  assign n10996 = n10994 & n10995 ;
  assign n10998 = n10996 ^ n10992 ;
  assign n10987 = n10813 ^ n10811 ;
  assign n10988 = n10814 ^ n10812 ;
  assign n10989 = n10987 & n10988 ;
  assign n10991 = n10989 ^ n10985 ;
  assign n11012 = n10998 ^ n10991 ;
  assign n10962 = n10809 ^ n10807 ;
  assign n10963 = n10810 ^ n10808 ;
  assign n10964 = n10962 & n10963 ;
  assign n10966 = n10964 ^ n10960 ;
  assign n10955 = n10805 ^ n10803 ;
  assign n10956 = n10806 ^ n10804 ;
  assign n10957 = n10955 & n10956 ;
  assign n10959 = n10957 ^ n10953 ;
  assign n10980 = n10966 ^ n10959 ;
  assign n11061 = n11012 ^ n10980 ;
  assign n10875 = n10801 ^ n10799 ;
  assign n10876 = n10802 ^ n10800 ;
  assign n10877 = n10875 & n10876 ;
  assign n10879 = n10877 ^ n10873 ;
  assign n10868 = n10797 ^ n10795 ;
  assign n10869 = n10798 ^ n10796 ;
  assign n10870 = n10868 & n10869 ;
  assign n10872 = n10870 ^ n10866 ;
  assign n10893 = n10879 ^ n10872 ;
  assign n10843 = n10793 ^ n10791 ;
  assign n10844 = n10794 ^ n10792 ;
  assign n10845 = n10843 & n10844 ;
  assign n10847 = n10845 ^ n10841 ;
  assign n10836 = n10789 ^ n10787 ;
  assign n10837 = n10790 ^ n10788 ;
  assign n10838 = n10836 & n10837 ;
  assign n10840 = n10838 ^ n10834 ;
  assign n10861 = n10847 ^ n10840 ;
  assign n10942 = n10893 ^ n10861 ;
  assign n11215 = n11061 ^ n10942 ;
  assign n11256 = n11239 ^ n11215 ;
  assign n11257 = n11256 ^ n10774 ;
  assign n9687 = n9510 ^ n9508 ;
  assign n9688 = n9511 ^ n9509 ;
  assign n9689 = n9687 & n9688 ;
  assign n9691 = n9689 ^ n9685 ;
  assign n9680 = n9506 ^ n9504 ;
  assign n9681 = n9507 ^ n9505 ;
  assign n9682 = n9680 & n9681 ;
  assign n9684 = n9682 ^ n9678 ;
  assign n9705 = n9691 ^ n9684 ;
  assign n9655 = n9502 ^ n9500 ;
  assign n9656 = n9503 ^ n9501 ;
  assign n9657 = n9655 & n9656 ;
  assign n9659 = n9657 ^ n9653 ;
  assign n9648 = n9498 ^ n9496 ;
  assign n9649 = n9499 ^ n9497 ;
  assign n9650 = n9648 & n9649 ;
  assign n9652 = n9650 ^ n9646 ;
  assign n9673 = n9659 ^ n9652 ;
  assign n9754 = n9705 ^ n9673 ;
  assign n9568 = n9494 ^ n9492 ;
  assign n9569 = n9495 ^ n9493 ;
  assign n9570 = n9568 & n9569 ;
  assign n9572 = n9570 ^ n9566 ;
  assign n9561 = n9490 ^ n9488 ;
  assign n9562 = n9491 ^ n9489 ;
  assign n9563 = n9561 & n9562 ;
  assign n9565 = n9563 ^ n9559 ;
  assign n9586 = n9572 ^ n9565 ;
  assign n9536 = n9486 ^ n9484 ;
  assign n9537 = n9487 ^ n9485 ;
  assign n9538 = n9536 & n9537 ;
  assign n9540 = n9538 ^ n9534 ;
  assign n9529 = n9482 ^ n9480 ;
  assign n9530 = n9483 ^ n9481 ;
  assign n9531 = n9529 & n9530 ;
  assign n9533 = n9531 ^ n9527 ;
  assign n9554 = n9540 ^ n9533 ;
  assign n9635 = n9586 ^ n9554 ;
  assign n9908 = n9754 ^ n9635 ;
  assign n9949 = n9932 ^ n9908 ;
  assign n9950 = n9949 ^ n9467 ;
  assign n12705 = n11257 ^ n9950 ;
  assign n12882 = n12801 ^ n12705 ;
  assign n12883 = n12882 ^ n8452 ;
  assign n11001 = n10817 ^ n10813 ;
  assign n11002 = n10818 ^ n10814 ;
  assign n11005 = n11001 & n11002 ;
  assign n10999 = n10815 ^ n10811 ;
  assign n11000 = n10816 ^ n10812 ;
  assign n11004 = n10999 & n11000 ;
  assign n11009 = n11005 ^ n11004 ;
  assign n11013 = n11011 ^ n11009 ;
  assign n11014 = n11013 ^ n10998 ;
  assign n10969 = n10809 ^ n10805 ;
  assign n10970 = n10810 ^ n10806 ;
  assign n10973 = n10969 & n10970 ;
  assign n10967 = n10807 ^ n10803 ;
  assign n10968 = n10808 ^ n10804 ;
  assign n10972 = n10967 & n10968 ;
  assign n10977 = n10973 ^ n10972 ;
  assign n10981 = n10979 ^ n10977 ;
  assign n10982 = n10981 ^ n10966 ;
  assign n11062 = n11014 ^ n10982 ;
  assign n10882 = n10801 ^ n10797 ;
  assign n10883 = n10802 ^ n10798 ;
  assign n10886 = n10882 & n10883 ;
  assign n10880 = n10799 ^ n10795 ;
  assign n10881 = n10800 ^ n10796 ;
  assign n10885 = n10880 & n10881 ;
  assign n10890 = n10886 ^ n10885 ;
  assign n10894 = n10892 ^ n10890 ;
  assign n10895 = n10894 ^ n10879 ;
  assign n10850 = n10793 ^ n10789 ;
  assign n10851 = n10794 ^ n10790 ;
  assign n10854 = n10850 & n10851 ;
  assign n10848 = n10791 ^ n10787 ;
  assign n10849 = n10792 ^ n10788 ;
  assign n10853 = n10848 & n10849 ;
  assign n10858 = n10854 ^ n10853 ;
  assign n10862 = n10860 ^ n10858 ;
  assign n10863 = n10862 ^ n10847 ;
  assign n10943 = n10895 ^ n10863 ;
  assign n11216 = n11062 ^ n10943 ;
  assign n11258 = n11240 ^ n11216 ;
  assign n11259 = n11258 ^ n10776 ;
  assign n9694 = n9510 ^ n9506 ;
  assign n9695 = n9511 ^ n9507 ;
  assign n9698 = n9694 & n9695 ;
  assign n9692 = n9508 ^ n9504 ;
  assign n9693 = n9509 ^ n9505 ;
  assign n9697 = n9692 & n9693 ;
  assign n9702 = n9698 ^ n9697 ;
  assign n9706 = n9704 ^ n9702 ;
  assign n9707 = n9706 ^ n9691 ;
  assign n9662 = n9502 ^ n9498 ;
  assign n9663 = n9503 ^ n9499 ;
  assign n9666 = n9662 & n9663 ;
  assign n9660 = n9500 ^ n9496 ;
  assign n9661 = n9501 ^ n9497 ;
  assign n9665 = n9660 & n9661 ;
  assign n9670 = n9666 ^ n9665 ;
  assign n9674 = n9672 ^ n9670 ;
  assign n9675 = n9674 ^ n9659 ;
  assign n9755 = n9707 ^ n9675 ;
  assign n9575 = n9494 ^ n9490 ;
  assign n9576 = n9495 ^ n9491 ;
  assign n9579 = n9575 & n9576 ;
  assign n9573 = n9492 ^ n9488 ;
  assign n9574 = n9493 ^ n9489 ;
  assign n9578 = n9573 & n9574 ;
  assign n9583 = n9579 ^ n9578 ;
  assign n9587 = n9585 ^ n9583 ;
  assign n9588 = n9587 ^ n9572 ;
  assign n9543 = n9486 ^ n9482 ;
  assign n9544 = n9487 ^ n9483 ;
  assign n9547 = n9543 & n9544 ;
  assign n9541 = n9484 ^ n9480 ;
  assign n9542 = n9485 ^ n9481 ;
  assign n9546 = n9541 & n9542 ;
  assign n9551 = n9547 ^ n9546 ;
  assign n9555 = n9553 ^ n9551 ;
  assign n9556 = n9555 ^ n9540 ;
  assign n9636 = n9588 ^ n9556 ;
  assign n9909 = n9755 ^ n9636 ;
  assign n9951 = n9933 ^ n9909 ;
  assign n9952 = n9951 ^ n9469 ;
  assign n12706 = n11259 ^ n9952 ;
  assign n12884 = n12802 ^ n12706 ;
  assign n12885 = n12884 ^ n8454 ;
  assign n11006 = n11001 ^ n10999 ;
  assign n11007 = n11002 ^ n11000 ;
  assign n11008 = n11006 & n11007 ;
  assign n11010 = n11008 ^ n11004 ;
  assign n11015 = n11012 ^ n11010 ;
  assign n11003 = n10998 ^ n10997 ;
  assign n11016 = n11015 ^ n11003 ;
  assign n10974 = n10969 ^ n10967 ;
  assign n10975 = n10970 ^ n10968 ;
  assign n10976 = n10974 & n10975 ;
  assign n10978 = n10976 ^ n10972 ;
  assign n10983 = n10980 ^ n10978 ;
  assign n10971 = n10966 ^ n10965 ;
  assign n10984 = n10983 ^ n10971 ;
  assign n11063 = n11016 ^ n10984 ;
  assign n10887 = n10882 ^ n10880 ;
  assign n10888 = n10883 ^ n10881 ;
  assign n10889 = n10887 & n10888 ;
  assign n10891 = n10889 ^ n10885 ;
  assign n10896 = n10893 ^ n10891 ;
  assign n10884 = n10879 ^ n10878 ;
  assign n10897 = n10896 ^ n10884 ;
  assign n10855 = n10850 ^ n10848 ;
  assign n10856 = n10851 ^ n10849 ;
  assign n10857 = n10855 & n10856 ;
  assign n10859 = n10857 ^ n10853 ;
  assign n10864 = n10861 ^ n10859 ;
  assign n10852 = n10847 ^ n10846 ;
  assign n10865 = n10864 ^ n10852 ;
  assign n10944 = n10897 ^ n10865 ;
  assign n11217 = n11063 ^ n10944 ;
  assign n11260 = n11241 ^ n11217 ;
  assign n11261 = n11260 ^ n10778 ;
  assign n9699 = n9694 ^ n9692 ;
  assign n9700 = n9695 ^ n9693 ;
  assign n9701 = n9699 & n9700 ;
  assign n9703 = n9701 ^ n9697 ;
  assign n9708 = n9705 ^ n9703 ;
  assign n9696 = n9691 ^ n9690 ;
  assign n9709 = n9708 ^ n9696 ;
  assign n9667 = n9662 ^ n9660 ;
  assign n9668 = n9663 ^ n9661 ;
  assign n9669 = n9667 & n9668 ;
  assign n9671 = n9669 ^ n9665 ;
  assign n9676 = n9673 ^ n9671 ;
  assign n9664 = n9659 ^ n9658 ;
  assign n9677 = n9676 ^ n9664 ;
  assign n9756 = n9709 ^ n9677 ;
  assign n9580 = n9575 ^ n9573 ;
  assign n9581 = n9576 ^ n9574 ;
  assign n9582 = n9580 & n9581 ;
  assign n9584 = n9582 ^ n9578 ;
  assign n9589 = n9586 ^ n9584 ;
  assign n9577 = n9572 ^ n9571 ;
  assign n9590 = n9589 ^ n9577 ;
  assign n9548 = n9543 ^ n9541 ;
  assign n9549 = n9544 ^ n9542 ;
  assign n9550 = n9548 & n9549 ;
  assign n9552 = n9550 ^ n9546 ;
  assign n9557 = n9554 ^ n9552 ;
  assign n9545 = n9540 ^ n9539 ;
  assign n9558 = n9557 ^ n9545 ;
  assign n9637 = n9590 ^ n9558 ;
  assign n9910 = n9756 ^ n9637 ;
  assign n9953 = n9934 ^ n9910 ;
  assign n9954 = n9953 ^ n9471 ;
  assign n12707 = n11261 ^ n9954 ;
  assign n12886 = n12803 ^ n12707 ;
  assign n12887 = n12886 ^ n8456 ;
  assign n11023 = n10817 ^ n10809 ;
  assign n11024 = n10818 ^ n10810 ;
  assign n11036 = n11023 & n11024 ;
  assign n11021 = n10815 ^ n10807 ;
  assign n11022 = n10816 ^ n10808 ;
  assign n11035 = n11021 & n11022 ;
  assign n11040 = n11036 ^ n11035 ;
  assign n11019 = n10813 ^ n10805 ;
  assign n11020 = n10814 ^ n10806 ;
  assign n11029 = n11019 & n11020 ;
  assign n11017 = n10811 ^ n10803 ;
  assign n11018 = n10812 ^ n10804 ;
  assign n11028 = n11017 & n11018 ;
  assign n11033 = n11029 ^ n11028 ;
  assign n11054 = n11040 ^ n11033 ;
  assign n11064 = n11060 ^ n11054 ;
  assign n11065 = n11064 ^ n11014 ;
  assign n10904 = n10801 ^ n10793 ;
  assign n10905 = n10802 ^ n10794 ;
  assign n10917 = n10904 & n10905 ;
  assign n10902 = n10799 ^ n10791 ;
  assign n10903 = n10800 ^ n10792 ;
  assign n10916 = n10902 & n10903 ;
  assign n10921 = n10917 ^ n10916 ;
  assign n10900 = n10797 ^ n10789 ;
  assign n10901 = n10798 ^ n10790 ;
  assign n10910 = n10900 & n10901 ;
  assign n10898 = n10795 ^ n10787 ;
  assign n10899 = n10796 ^ n10788 ;
  assign n10909 = n10898 & n10899 ;
  assign n10914 = n10910 ^ n10909 ;
  assign n10935 = n10921 ^ n10914 ;
  assign n10945 = n10941 ^ n10935 ;
  assign n10946 = n10945 ^ n10895 ;
  assign n11218 = n11065 ^ n10946 ;
  assign n11262 = n11242 ^ n11218 ;
  assign n11263 = n11262 ^ n10780 ;
  assign n9716 = n9510 ^ n9502 ;
  assign n9717 = n9511 ^ n9503 ;
  assign n9729 = n9716 & n9717 ;
  assign n9714 = n9508 ^ n9500 ;
  assign n9715 = n9509 ^ n9501 ;
  assign n9728 = n9714 & n9715 ;
  assign n9733 = n9729 ^ n9728 ;
  assign n9712 = n9506 ^ n9498 ;
  assign n9713 = n9507 ^ n9499 ;
  assign n9722 = n9712 & n9713 ;
  assign n9710 = n9504 ^ n9496 ;
  assign n9711 = n9505 ^ n9497 ;
  assign n9721 = n9710 & n9711 ;
  assign n9726 = n9722 ^ n9721 ;
  assign n9747 = n9733 ^ n9726 ;
  assign n9757 = n9753 ^ n9747 ;
  assign n9758 = n9757 ^ n9707 ;
  assign n9597 = n9494 ^ n9486 ;
  assign n9598 = n9495 ^ n9487 ;
  assign n9610 = n9597 & n9598 ;
  assign n9595 = n9492 ^ n9484 ;
  assign n9596 = n9493 ^ n9485 ;
  assign n9609 = n9595 & n9596 ;
  assign n9614 = n9610 ^ n9609 ;
  assign n9593 = n9490 ^ n9482 ;
  assign n9594 = n9491 ^ n9483 ;
  assign n9603 = n9593 & n9594 ;
  assign n9591 = n9488 ^ n9480 ;
  assign n9592 = n9489 ^ n9481 ;
  assign n9602 = n9591 & n9592 ;
  assign n9607 = n9603 ^ n9602 ;
  assign n9628 = n9614 ^ n9607 ;
  assign n9638 = n9634 ^ n9628 ;
  assign n9639 = n9638 ^ n9588 ;
  assign n9911 = n9758 ^ n9639 ;
  assign n9955 = n9935 ^ n9911 ;
  assign n9956 = n9955 ^ n9473 ;
  assign n12708 = n11263 ^ n9956 ;
  assign n12888 = n12804 ^ n12708 ;
  assign n12889 = n12888 ^ n8458 ;
  assign n11037 = n11023 ^ n11021 ;
  assign n11038 = n11024 ^ n11022 ;
  assign n11039 = n11037 & n11038 ;
  assign n11041 = n11039 ^ n11035 ;
  assign n11030 = n11019 ^ n11017 ;
  assign n11031 = n11020 ^ n11018 ;
  assign n11032 = n11030 & n11031 ;
  assign n11034 = n11032 ^ n11028 ;
  assign n11055 = n11041 ^ n11034 ;
  assign n11066 = n11061 ^ n11055 ;
  assign n11067 = n11066 ^ n11016 ;
  assign n10918 = n10904 ^ n10902 ;
  assign n10919 = n10905 ^ n10903 ;
  assign n10920 = n10918 & n10919 ;
  assign n10922 = n10920 ^ n10916 ;
  assign n10911 = n10900 ^ n10898 ;
  assign n10912 = n10901 ^ n10899 ;
  assign n10913 = n10911 & n10912 ;
  assign n10915 = n10913 ^ n10909 ;
  assign n10936 = n10922 ^ n10915 ;
  assign n10947 = n10942 ^ n10936 ;
  assign n10948 = n10947 ^ n10897 ;
  assign n11219 = n11067 ^ n10948 ;
  assign n11264 = n11243 ^ n11219 ;
  assign n11265 = n11264 ^ n10782 ;
  assign n9730 = n9716 ^ n9714 ;
  assign n9731 = n9717 ^ n9715 ;
  assign n9732 = n9730 & n9731 ;
  assign n9734 = n9732 ^ n9728 ;
  assign n9723 = n9712 ^ n9710 ;
  assign n9724 = n9713 ^ n9711 ;
  assign n9725 = n9723 & n9724 ;
  assign n9727 = n9725 ^ n9721 ;
  assign n9748 = n9734 ^ n9727 ;
  assign n9759 = n9754 ^ n9748 ;
  assign n9760 = n9759 ^ n9709 ;
  assign n9611 = n9597 ^ n9595 ;
  assign n9612 = n9598 ^ n9596 ;
  assign n9613 = n9611 & n9612 ;
  assign n9615 = n9613 ^ n9609 ;
  assign n9604 = n9593 ^ n9591 ;
  assign n9605 = n9594 ^ n9592 ;
  assign n9606 = n9604 & n9605 ;
  assign n9608 = n9606 ^ n9602 ;
  assign n9629 = n9615 ^ n9608 ;
  assign n9640 = n9635 ^ n9629 ;
  assign n9641 = n9640 ^ n9590 ;
  assign n9912 = n9760 ^ n9641 ;
  assign n9957 = n9936 ^ n9912 ;
  assign n9958 = n9957 ^ n9475 ;
  assign n12709 = n11265 ^ n9958 ;
  assign n12890 = n12805 ^ n12709 ;
  assign n12891 = n12890 ^ n8460 ;
  assign n11044 = n11023 ^ n11019 ;
  assign n11045 = n11024 ^ n11020 ;
  assign n11048 = n11044 & n11045 ;
  assign n11042 = n11021 ^ n11017 ;
  assign n11043 = n11022 ^ n11018 ;
  assign n11047 = n11042 & n11043 ;
  assign n11052 = n11048 ^ n11047 ;
  assign n11056 = n11054 ^ n11052 ;
  assign n11057 = n11056 ^ n11041 ;
  assign n11068 = n11062 ^ n11057 ;
  assign n11026 = n11016 ^ n11011 ;
  assign n11069 = n11068 ^ n11026 ;
  assign n10925 = n10904 ^ n10900 ;
  assign n10926 = n10905 ^ n10901 ;
  assign n10929 = n10925 & n10926 ;
  assign n10923 = n10902 ^ n10898 ;
  assign n10924 = n10903 ^ n10899 ;
  assign n10928 = n10923 & n10924 ;
  assign n10933 = n10929 ^ n10928 ;
  assign n10937 = n10935 ^ n10933 ;
  assign n10938 = n10937 ^ n10922 ;
  assign n10949 = n10943 ^ n10938 ;
  assign n10907 = n10897 ^ n10892 ;
  assign n10950 = n10949 ^ n10907 ;
  assign n11220 = n11069 ^ n10950 ;
  assign n11266 = n11244 ^ n11220 ;
  assign n11267 = n11266 ^ n10784 ;
  assign n9737 = n9716 ^ n9712 ;
  assign n9738 = n9717 ^ n9713 ;
  assign n9741 = n9737 & n9738 ;
  assign n9735 = n9714 ^ n9710 ;
  assign n9736 = n9715 ^ n9711 ;
  assign n9740 = n9735 & n9736 ;
  assign n9745 = n9741 ^ n9740 ;
  assign n9749 = n9747 ^ n9745 ;
  assign n9750 = n9749 ^ n9734 ;
  assign n9761 = n9755 ^ n9750 ;
  assign n9719 = n9709 ^ n9704 ;
  assign n9762 = n9761 ^ n9719 ;
  assign n9618 = n9597 ^ n9593 ;
  assign n9619 = n9598 ^ n9594 ;
  assign n9622 = n9618 & n9619 ;
  assign n9616 = n9595 ^ n9591 ;
  assign n9617 = n9596 ^ n9592 ;
  assign n9621 = n9616 & n9617 ;
  assign n9626 = n9622 ^ n9621 ;
  assign n9630 = n9628 ^ n9626 ;
  assign n9631 = n9630 ^ n9615 ;
  assign n9642 = n9636 ^ n9631 ;
  assign n9600 = n9590 ^ n9585 ;
  assign n9643 = n9642 ^ n9600 ;
  assign n9913 = n9762 ^ n9643 ;
  assign n9959 = n9937 ^ n9913 ;
  assign n9960 = n9959 ^ n9477 ;
  assign n12710 = n11267 ^ n9960 ;
  assign n12892 = n12806 ^ n12710 ;
  assign n12893 = n12892 ^ n8462 ;
  assign n11049 = n11044 ^ n11042 ;
  assign n11050 = n11045 ^ n11043 ;
  assign n11051 = n11049 & n11050 ;
  assign n11053 = n11051 ^ n11047 ;
  assign n11058 = n11055 ^ n11053 ;
  assign n11046 = n11041 ^ n11040 ;
  assign n11059 = n11058 ^ n11046 ;
  assign n11070 = n11063 ^ n11059 ;
  assign n11025 = n11016 ^ n11014 ;
  assign n11027 = n11025 ^ n11012 ;
  assign n11071 = n11070 ^ n11027 ;
  assign n10930 = n10925 ^ n10923 ;
  assign n10931 = n10926 ^ n10924 ;
  assign n10932 = n10930 & n10931 ;
  assign n10934 = n10932 ^ n10928 ;
  assign n10939 = n10936 ^ n10934 ;
  assign n10927 = n10922 ^ n10921 ;
  assign n10940 = n10939 ^ n10927 ;
  assign n10951 = n10944 ^ n10940 ;
  assign n10906 = n10897 ^ n10895 ;
  assign n10908 = n10906 ^ n10893 ;
  assign n10952 = n10951 ^ n10908 ;
  assign n11221 = n11071 ^ n10952 ;
  assign n11268 = n11245 ^ n11221 ;
  assign n11269 = n11268 ^ n10786 ;
  assign n9742 = n9737 ^ n9735 ;
  assign n9743 = n9738 ^ n9736 ;
  assign n9744 = n9742 & n9743 ;
  assign n9746 = n9744 ^ n9740 ;
  assign n9751 = n9748 ^ n9746 ;
  assign n9739 = n9734 ^ n9733 ;
  assign n9752 = n9751 ^ n9739 ;
  assign n9763 = n9756 ^ n9752 ;
  assign n9718 = n9709 ^ n9707 ;
  assign n9720 = n9718 ^ n9705 ;
  assign n9764 = n9763 ^ n9720 ;
  assign n9623 = n9618 ^ n9616 ;
  assign n9624 = n9619 ^ n9617 ;
  assign n9625 = n9623 & n9624 ;
  assign n9627 = n9625 ^ n9621 ;
  assign n9632 = n9629 ^ n9627 ;
  assign n9620 = n9615 ^ n9614 ;
  assign n9633 = n9632 ^ n9620 ;
  assign n9644 = n9637 ^ n9633 ;
  assign n9599 = n9590 ^ n9588 ;
  assign n9601 = n9599 ^ n9586 ;
  assign n9645 = n9644 ^ n9601 ;
  assign n9914 = n9764 ^ n9645 ;
  assign n9961 = n9938 ^ n9914 ;
  assign n9962 = n9961 ^ n9479 ;
  assign n12711 = n11269 ^ n9962 ;
  assign n12894 = n12807 ^ n12711 ;
  assign n12895 = n12894 ^ n8464 ;
  assign n11086 = n10817 ^ n10801 ;
  assign n11087 = n10818 ^ n10802 ;
  assign n11135 = n11086 & n11087 ;
  assign n11084 = n10815 ^ n10799 ;
  assign n11085 = n10816 ^ n10800 ;
  assign n11134 = n11084 & n11085 ;
  assign n11139 = n11135 ^ n11134 ;
  assign n11082 = n10813 ^ n10797 ;
  assign n11083 = n10814 ^ n10798 ;
  assign n11128 = n11082 & n11083 ;
  assign n11080 = n10811 ^ n10795 ;
  assign n11081 = n10812 ^ n10796 ;
  assign n11127 = n11080 & n11081 ;
  assign n11132 = n11128 ^ n11127 ;
  assign n11153 = n11139 ^ n11132 ;
  assign n11078 = n10809 ^ n10793 ;
  assign n11079 = n10810 ^ n10794 ;
  assign n11103 = n11078 & n11079 ;
  assign n11076 = n10807 ^ n10791 ;
  assign n11077 = n10808 ^ n10792 ;
  assign n11102 = n11076 & n11077 ;
  assign n11107 = n11103 ^ n11102 ;
  assign n11074 = n10805 ^ n10789 ;
  assign n11075 = n10806 ^ n10790 ;
  assign n11096 = n11074 & n11075 ;
  assign n11072 = n10803 ^ n10787 ;
  assign n11073 = n10804 ^ n10788 ;
  assign n11095 = n11072 & n11073 ;
  assign n11100 = n11096 ^ n11095 ;
  assign n11121 = n11107 ^ n11100 ;
  assign n11202 = n11153 ^ n11121 ;
  assign n11222 = n11214 ^ n11202 ;
  assign n11223 = n11222 ^ n11065 ;
  assign n11270 = n11246 ^ n11223 ;
  assign n10826 = n10780 ^ n10763 ;
  assign n11271 = n11270 ^ n10826 ;
  assign n9779 = n9510 ^ n9494 ;
  assign n9780 = n9511 ^ n9495 ;
  assign n9828 = n9779 & n9780 ;
  assign n9777 = n9508 ^ n9492 ;
  assign n9778 = n9509 ^ n9493 ;
  assign n9827 = n9777 & n9778 ;
  assign n9832 = n9828 ^ n9827 ;
  assign n9775 = n9506 ^ n9490 ;
  assign n9776 = n9507 ^ n9491 ;
  assign n9821 = n9775 & n9776 ;
  assign n9773 = n9504 ^ n9488 ;
  assign n9774 = n9505 ^ n9489 ;
  assign n9820 = n9773 & n9774 ;
  assign n9825 = n9821 ^ n9820 ;
  assign n9846 = n9832 ^ n9825 ;
  assign n9771 = n9502 ^ n9486 ;
  assign n9772 = n9503 ^ n9487 ;
  assign n9796 = n9771 & n9772 ;
  assign n9769 = n9500 ^ n9484 ;
  assign n9770 = n9501 ^ n9485 ;
  assign n9795 = n9769 & n9770 ;
  assign n9800 = n9796 ^ n9795 ;
  assign n9767 = n9498 ^ n9482 ;
  assign n9768 = n9499 ^ n9483 ;
  assign n9789 = n9767 & n9768 ;
  assign n9765 = n9496 ^ n9480 ;
  assign n9766 = n9497 ^ n9481 ;
  assign n9788 = n9765 & n9766 ;
  assign n9793 = n9789 ^ n9788 ;
  assign n9814 = n9800 ^ n9793 ;
  assign n9895 = n9846 ^ n9814 ;
  assign n9915 = n9907 ^ n9895 ;
  assign n9916 = n9915 ^ n9758 ;
  assign n9963 = n9939 ^ n9916 ;
  assign n9519 = n9473 ^ n9456 ;
  assign n9964 = n9963 ^ n9519 ;
  assign n12712 = n11271 ^ n9964 ;
  assign n12896 = n12808 ^ n12712 ;
  assign n12897 = n12896 ^ n8466 ;
  assign n11136 = n11086 ^ n11084 ;
  assign n11137 = n11087 ^ n11085 ;
  assign n11138 = n11136 & n11137 ;
  assign n11140 = n11138 ^ n11134 ;
  assign n11129 = n11082 ^ n11080 ;
  assign n11130 = n11083 ^ n11081 ;
  assign n11131 = n11129 & n11130 ;
  assign n11133 = n11131 ^ n11127 ;
  assign n11154 = n11140 ^ n11133 ;
  assign n11104 = n11078 ^ n11076 ;
  assign n11105 = n11079 ^ n11077 ;
  assign n11106 = n11104 & n11105 ;
  assign n11108 = n11106 ^ n11102 ;
  assign n11097 = n11074 ^ n11072 ;
  assign n11098 = n11075 ^ n11073 ;
  assign n11099 = n11097 & n11098 ;
  assign n11101 = n11099 ^ n11095 ;
  assign n11122 = n11108 ^ n11101 ;
  assign n11203 = n11154 ^ n11122 ;
  assign n11224 = n11215 ^ n11203 ;
  assign n11225 = n11224 ^ n11067 ;
  assign n11272 = n11247 ^ n11225 ;
  assign n10827 = n10782 ^ n10764 ;
  assign n11273 = n11272 ^ n10827 ;
  assign n9829 = n9779 ^ n9777 ;
  assign n9830 = n9780 ^ n9778 ;
  assign n9831 = n9829 & n9830 ;
  assign n9833 = n9831 ^ n9827 ;
  assign n9822 = n9775 ^ n9773 ;
  assign n9823 = n9776 ^ n9774 ;
  assign n9824 = n9822 & n9823 ;
  assign n9826 = n9824 ^ n9820 ;
  assign n9847 = n9833 ^ n9826 ;
  assign n9797 = n9771 ^ n9769 ;
  assign n9798 = n9772 ^ n9770 ;
  assign n9799 = n9797 & n9798 ;
  assign n9801 = n9799 ^ n9795 ;
  assign n9790 = n9767 ^ n9765 ;
  assign n9791 = n9768 ^ n9766 ;
  assign n9792 = n9790 & n9791 ;
  assign n9794 = n9792 ^ n9788 ;
  assign n9815 = n9801 ^ n9794 ;
  assign n9896 = n9847 ^ n9815 ;
  assign n9917 = n9908 ^ n9896 ;
  assign n9918 = n9917 ^ n9760 ;
  assign n9965 = n9940 ^ n9918 ;
  assign n9520 = n9475 ^ n9457 ;
  assign n9966 = n9965 ^ n9520 ;
  assign n12713 = n11273 ^ n9966 ;
  assign n12898 = n12809 ^ n12713 ;
  assign n12899 = n12898 ^ n8468 ;
  assign n11143 = n11086 ^ n11082 ;
  assign n11144 = n11087 ^ n11083 ;
  assign n11147 = n11143 & n11144 ;
  assign n11141 = n11084 ^ n11080 ;
  assign n11142 = n11085 ^ n11081 ;
  assign n11146 = n11141 & n11142 ;
  assign n11151 = n11147 ^ n11146 ;
  assign n11155 = n11153 ^ n11151 ;
  assign n11156 = n11155 ^ n11140 ;
  assign n11111 = n11078 ^ n11074 ;
  assign n11112 = n11079 ^ n11075 ;
  assign n11115 = n11111 & n11112 ;
  assign n11109 = n11076 ^ n11072 ;
  assign n11110 = n11077 ^ n11073 ;
  assign n11114 = n11109 & n11110 ;
  assign n11119 = n11115 ^ n11114 ;
  assign n11123 = n11121 ^ n11119 ;
  assign n11124 = n11123 ^ n11108 ;
  assign n11204 = n11156 ^ n11124 ;
  assign n11226 = n11216 ^ n11204 ;
  assign n11227 = n11226 ^ n11069 ;
  assign n11274 = n11248 ^ n11227 ;
  assign n10828 = n10784 ^ n10765 ;
  assign n11275 = n11274 ^ n10828 ;
  assign n9836 = n9779 ^ n9775 ;
  assign n9837 = n9780 ^ n9776 ;
  assign n9840 = n9836 & n9837 ;
  assign n9834 = n9777 ^ n9773 ;
  assign n9835 = n9778 ^ n9774 ;
  assign n9839 = n9834 & n9835 ;
  assign n9844 = n9840 ^ n9839 ;
  assign n9848 = n9846 ^ n9844 ;
  assign n9849 = n9848 ^ n9833 ;
  assign n9804 = n9771 ^ n9767 ;
  assign n9805 = n9772 ^ n9768 ;
  assign n9808 = n9804 & n9805 ;
  assign n9802 = n9769 ^ n9765 ;
  assign n9803 = n9770 ^ n9766 ;
  assign n9807 = n9802 & n9803 ;
  assign n9812 = n9808 ^ n9807 ;
  assign n9816 = n9814 ^ n9812 ;
  assign n9817 = n9816 ^ n9801 ;
  assign n9897 = n9849 ^ n9817 ;
  assign n9919 = n9909 ^ n9897 ;
  assign n9920 = n9919 ^ n9762 ;
  assign n9967 = n9941 ^ n9920 ;
  assign n9521 = n9477 ^ n9458 ;
  assign n9968 = n9967 ^ n9521 ;
  assign n12714 = n11275 ^ n9968 ;
  assign n12900 = n12810 ^ n12714 ;
  assign n12901 = n12900 ^ n8470 ;
  assign n11148 = n11143 ^ n11141 ;
  assign n11149 = n11144 ^ n11142 ;
  assign n11150 = n11148 & n11149 ;
  assign n11152 = n11150 ^ n11146 ;
  assign n11157 = n11154 ^ n11152 ;
  assign n11145 = n11140 ^ n11139 ;
  assign n11158 = n11157 ^ n11145 ;
  assign n11116 = n11111 ^ n11109 ;
  assign n11117 = n11112 ^ n11110 ;
  assign n11118 = n11116 & n11117 ;
  assign n11120 = n11118 ^ n11114 ;
  assign n11125 = n11122 ^ n11120 ;
  assign n11113 = n11108 ^ n11107 ;
  assign n11126 = n11125 ^ n11113 ;
  assign n11205 = n11158 ^ n11126 ;
  assign n11228 = n11217 ^ n11205 ;
  assign n11229 = n11228 ^ n11071 ;
  assign n11276 = n11249 ^ n11229 ;
  assign n10829 = n10786 ^ n10766 ;
  assign n11277 = n11276 ^ n10829 ;
  assign n9841 = n9836 ^ n9834 ;
  assign n9842 = n9837 ^ n9835 ;
  assign n9843 = n9841 & n9842 ;
  assign n9845 = n9843 ^ n9839 ;
  assign n9850 = n9847 ^ n9845 ;
  assign n9838 = n9833 ^ n9832 ;
  assign n9851 = n9850 ^ n9838 ;
  assign n9809 = n9804 ^ n9802 ;
  assign n9810 = n9805 ^ n9803 ;
  assign n9811 = n9809 & n9810 ;
  assign n9813 = n9811 ^ n9807 ;
  assign n9818 = n9815 ^ n9813 ;
  assign n9806 = n9801 ^ n9800 ;
  assign n9819 = n9818 ^ n9806 ;
  assign n9898 = n9851 ^ n9819 ;
  assign n9921 = n9910 ^ n9898 ;
  assign n9922 = n9921 ^ n9764 ;
  assign n9969 = n9942 ^ n9922 ;
  assign n9522 = n9479 ^ n9459 ;
  assign n9970 = n9969 ^ n9522 ;
  assign n12715 = n11277 ^ n9970 ;
  assign n12902 = n12811 ^ n12715 ;
  assign n12903 = n12902 ^ n8472 ;
  assign n11165 = n11086 ^ n11078 ;
  assign n11166 = n11087 ^ n11079 ;
  assign n11178 = n11165 & n11166 ;
  assign n11163 = n11084 ^ n11076 ;
  assign n11164 = n11085 ^ n11077 ;
  assign n11177 = n11163 & n11164 ;
  assign n11182 = n11178 ^ n11177 ;
  assign n11161 = n11082 ^ n11074 ;
  assign n11162 = n11083 ^ n11075 ;
  assign n11171 = n11161 & n11162 ;
  assign n11159 = n11080 ^ n11072 ;
  assign n11160 = n11081 ^ n11073 ;
  assign n11170 = n11159 & n11160 ;
  assign n11175 = n11171 ^ n11170 ;
  assign n11196 = n11182 ^ n11175 ;
  assign n11206 = n11202 ^ n11196 ;
  assign n11207 = n11206 ^ n11156 ;
  assign n11230 = n11218 ^ n11207 ;
  assign n11091 = n11069 ^ n11060 ;
  assign n11231 = n11230 ^ n11091 ;
  assign n11278 = n11250 ^ n11231 ;
  assign n10822 = n10784 ^ n10772 ;
  assign n10830 = n10822 ^ n10767 ;
  assign n11279 = n11278 ^ n10830 ;
  assign n9858 = n9779 ^ n9771 ;
  assign n9859 = n9780 ^ n9772 ;
  assign n9871 = n9858 & n9859 ;
  assign n9856 = n9777 ^ n9769 ;
  assign n9857 = n9778 ^ n9770 ;
  assign n9870 = n9856 & n9857 ;
  assign n9875 = n9871 ^ n9870 ;
  assign n9854 = n9775 ^ n9767 ;
  assign n9855 = n9776 ^ n9768 ;
  assign n9864 = n9854 & n9855 ;
  assign n9852 = n9773 ^ n9765 ;
  assign n9853 = n9774 ^ n9766 ;
  assign n9863 = n9852 & n9853 ;
  assign n9868 = n9864 ^ n9863 ;
  assign n9889 = n9875 ^ n9868 ;
  assign n9899 = n9895 ^ n9889 ;
  assign n9900 = n9899 ^ n9849 ;
  assign n9923 = n9911 ^ n9900 ;
  assign n9784 = n9762 ^ n9753 ;
  assign n9924 = n9923 ^ n9784 ;
  assign n9971 = n9943 ^ n9924 ;
  assign n9515 = n9477 ^ n9465 ;
  assign n9523 = n9515 ^ n9460 ;
  assign n9972 = n9971 ^ n9523 ;
  assign n12716 = n11279 ^ n9972 ;
  assign n12904 = n12812 ^ n12716 ;
  assign n12905 = n12904 ^ n8474 ;
  assign n11179 = n11165 ^ n11163 ;
  assign n11180 = n11166 ^ n11164 ;
  assign n11181 = n11179 & n11180 ;
  assign n11183 = n11181 ^ n11177 ;
  assign n11172 = n11161 ^ n11159 ;
  assign n11173 = n11162 ^ n11160 ;
  assign n11174 = n11172 & n11173 ;
  assign n11176 = n11174 ^ n11170 ;
  assign n11197 = n11183 ^ n11176 ;
  assign n11208 = n11203 ^ n11197 ;
  assign n11209 = n11208 ^ n11158 ;
  assign n11232 = n11219 ^ n11209 ;
  assign n11092 = n11071 ^ n11061 ;
  assign n11233 = n11232 ^ n11092 ;
  assign n11280 = n11251 ^ n11233 ;
  assign n10823 = n10786 ^ n10774 ;
  assign n10831 = n10823 ^ n10768 ;
  assign n11281 = n11280 ^ n10831 ;
  assign n9872 = n9858 ^ n9856 ;
  assign n9873 = n9859 ^ n9857 ;
  assign n9874 = n9872 & n9873 ;
  assign n9876 = n9874 ^ n9870 ;
  assign n9865 = n9854 ^ n9852 ;
  assign n9866 = n9855 ^ n9853 ;
  assign n9867 = n9865 & n9866 ;
  assign n9869 = n9867 ^ n9863 ;
  assign n9890 = n9876 ^ n9869 ;
  assign n9901 = n9896 ^ n9890 ;
  assign n9902 = n9901 ^ n9851 ;
  assign n9925 = n9912 ^ n9902 ;
  assign n9785 = n9764 ^ n9754 ;
  assign n9926 = n9925 ^ n9785 ;
  assign n9973 = n9944 ^ n9926 ;
  assign n9516 = n9479 ^ n9467 ;
  assign n9524 = n9516 ^ n9461 ;
  assign n9974 = n9973 ^ n9524 ;
  assign n12717 = n11281 ^ n9974 ;
  assign n12906 = n12813 ^ n12717 ;
  assign n12907 = n12906 ^ n8476 ;
  assign n11186 = n11165 ^ n11161 ;
  assign n11187 = n11166 ^ n11162 ;
  assign n11190 = n11186 & n11187 ;
  assign n11184 = n11163 ^ n11159 ;
  assign n11185 = n11164 ^ n11160 ;
  assign n11189 = n11184 & n11185 ;
  assign n11194 = n11190 ^ n11189 ;
  assign n11198 = n11196 ^ n11194 ;
  assign n11199 = n11198 ^ n11183 ;
  assign n11210 = n11204 ^ n11199 ;
  assign n11168 = n11158 ^ n11153 ;
  assign n11211 = n11210 ^ n11168 ;
  assign n11234 = n11220 ^ n11211 ;
  assign n11089 = n11071 ^ n11065 ;
  assign n11093 = n11089 ^ n11062 ;
  assign n11235 = n11234 ^ n11093 ;
  assign n11282 = n11252 ^ n11235 ;
  assign n10820 = n10786 ^ n10780 ;
  assign n10824 = n10820 ^ n10776 ;
  assign n10832 = n10824 ^ n10769 ;
  assign n11283 = n11282 ^ n10832 ;
  assign n9879 = n9858 ^ n9854 ;
  assign n9880 = n9859 ^ n9855 ;
  assign n9883 = n9879 & n9880 ;
  assign n9877 = n9856 ^ n9852 ;
  assign n9878 = n9857 ^ n9853 ;
  assign n9882 = n9877 & n9878 ;
  assign n9887 = n9883 ^ n9882 ;
  assign n9891 = n9889 ^ n9887 ;
  assign n9892 = n9891 ^ n9876 ;
  assign n9903 = n9897 ^ n9892 ;
  assign n9861 = n9851 ^ n9846 ;
  assign n9904 = n9903 ^ n9861 ;
  assign n9927 = n9913 ^ n9904 ;
  assign n9782 = n9764 ^ n9758 ;
  assign n9786 = n9782 ^ n9755 ;
  assign n9928 = n9927 ^ n9786 ;
  assign n9975 = n9945 ^ n9928 ;
  assign n9513 = n9479 ^ n9473 ;
  assign n9517 = n9513 ^ n9469 ;
  assign n9525 = n9517 ^ n9462 ;
  assign n9976 = n9975 ^ n9525 ;
  assign n12718 = n11283 ^ n9976 ;
  assign n12908 = n12814 ^ n12718 ;
  assign n12909 = n12908 ^ n8478 ;
  assign n11191 = n11186 ^ n11184 ;
  assign n11192 = n11187 ^ n11185 ;
  assign n11193 = n11191 & n11192 ;
  assign n11195 = n11193 ^ n11189 ;
  assign n11200 = n11197 ^ n11195 ;
  assign n11188 = n11183 ^ n11182 ;
  assign n11201 = n11200 ^ n11188 ;
  assign n11212 = n11205 ^ n11201 ;
  assign n11167 = n11158 ^ n11156 ;
  assign n11169 = n11167 ^ n11154 ;
  assign n11213 = n11212 ^ n11169 ;
  assign n11236 = n11221 ^ n11213 ;
  assign n11088 = n11071 ^ n11069 ;
  assign n11090 = n11088 ^ n11067 ;
  assign n11094 = n11090 ^ n11063 ;
  assign n11237 = n11236 ^ n11094 ;
  assign n11284 = n11253 ^ n11237 ;
  assign n10819 = n10786 ^ n10784 ;
  assign n10821 = n10819 ^ n10782 ;
  assign n10825 = n10821 ^ n10778 ;
  assign n10833 = n10825 ^ n10770 ;
  assign n11285 = n11284 ^ n10833 ;
  assign n9884 = n9879 ^ n9877 ;
  assign n9885 = n9880 ^ n9878 ;
  assign n9886 = n9884 & n9885 ;
  assign n9888 = n9886 ^ n9882 ;
  assign n9893 = n9890 ^ n9888 ;
  assign n9881 = n9876 ^ n9875 ;
  assign n9894 = n9893 ^ n9881 ;
  assign n9905 = n9898 ^ n9894 ;
  assign n9860 = n9851 ^ n9849 ;
  assign n9862 = n9860 ^ n9847 ;
  assign n9906 = n9905 ^ n9862 ;
  assign n9929 = n9914 ^ n9906 ;
  assign n9781 = n9764 ^ n9762 ;
  assign n9783 = n9781 ^ n9760 ;
  assign n9787 = n9783 ^ n9756 ;
  assign n9930 = n9929 ^ n9787 ;
  assign n9977 = n9946 ^ n9930 ;
  assign n9512 = n9479 ^ n9477 ;
  assign n9514 = n9512 ^ n9475 ;
  assign n9518 = n9514 ^ n9471 ;
  assign n9526 = n9518 ^ n9463 ;
  assign n9978 = n9977 ^ n9526 ;
  assign n12719 = n11285 ^ n9978 ;
  assign n12910 = n12815 ^ n12719 ;
  assign n12911 = n12910 ^ n8480 ;
  assign n11348 = n8607 ^ n8543 ;
  assign n11349 = n8608 ^ n8544 ;
  assign n11944 = n11348 & n11349 ;
  assign n11346 = n8605 ^ n8541 ;
  assign n11347 = n8606 ^ n8542 ;
  assign n11943 = n11346 & n11347 ;
  assign n11948 = n11944 ^ n11943 ;
  assign n11344 = n8603 ^ n8539 ;
  assign n11345 = n8604 ^ n8540 ;
  assign n11937 = n11344 & n11345 ;
  assign n11342 = n8601 ^ n8537 ;
  assign n11343 = n8602 ^ n8538 ;
  assign n11936 = n11342 & n11343 ;
  assign n11941 = n11937 ^ n11936 ;
  assign n11962 = n11948 ^ n11941 ;
  assign n11340 = n8599 ^ n8535 ;
  assign n11341 = n8600 ^ n8536 ;
  assign n11912 = n11340 & n11341 ;
  assign n11338 = n8597 ^ n8533 ;
  assign n11339 = n8598 ^ n8534 ;
  assign n11911 = n11338 & n11339 ;
  assign n11916 = n11912 ^ n11911 ;
  assign n11336 = n8595 ^ n8531 ;
  assign n11337 = n8596 ^ n8532 ;
  assign n11905 = n11336 & n11337 ;
  assign n11334 = n8593 ^ n8529 ;
  assign n11335 = n8594 ^ n8530 ;
  assign n11904 = n11334 & n11335 ;
  assign n11909 = n11905 ^ n11904 ;
  assign n11930 = n11916 ^ n11909 ;
  assign n12011 = n11962 ^ n11930 ;
  assign n11332 = n8591 ^ n8527 ;
  assign n11333 = n8592 ^ n8528 ;
  assign n11825 = n11332 & n11333 ;
  assign n11330 = n8589 ^ n8525 ;
  assign n11331 = n8590 ^ n8526 ;
  assign n11824 = n11330 & n11331 ;
  assign n11829 = n11825 ^ n11824 ;
  assign n11328 = n8587 ^ n8523 ;
  assign n11329 = n8588 ^ n8524 ;
  assign n11818 = n11328 & n11329 ;
  assign n11326 = n8585 ^ n8521 ;
  assign n11327 = n8586 ^ n8522 ;
  assign n11817 = n11326 & n11327 ;
  assign n11822 = n11818 ^ n11817 ;
  assign n11843 = n11829 ^ n11822 ;
  assign n11324 = n8583 ^ n8519 ;
  assign n11325 = n8584 ^ n8520 ;
  assign n11793 = n11324 & n11325 ;
  assign n11322 = n8581 ^ n8517 ;
  assign n11323 = n8582 ^ n8518 ;
  assign n11792 = n11322 & n11323 ;
  assign n11797 = n11793 ^ n11792 ;
  assign n11320 = n8579 ^ n8515 ;
  assign n11321 = n8580 ^ n8516 ;
  assign n11786 = n11320 & n11321 ;
  assign n11318 = n8577 ^ n8513 ;
  assign n11319 = n8578 ^ n8514 ;
  assign n11785 = n11318 & n11319 ;
  assign n11790 = n11786 ^ n11785 ;
  assign n11811 = n11797 ^ n11790 ;
  assign n11892 = n11843 ^ n11811 ;
  assign n12165 = n12011 ^ n11892 ;
  assign n11316 = n8575 ^ n8511 ;
  assign n11317 = n8576 ^ n8512 ;
  assign n11540 = n11316 & n11317 ;
  assign n11314 = n8573 ^ n8509 ;
  assign n11315 = n8574 ^ n8510 ;
  assign n11539 = n11314 & n11315 ;
  assign n11544 = n11540 ^ n11539 ;
  assign n11312 = n8571 ^ n8507 ;
  assign n11313 = n8572 ^ n8508 ;
  assign n11533 = n11312 & n11313 ;
  assign n11310 = n8569 ^ n8505 ;
  assign n11311 = n8570 ^ n8506 ;
  assign n11532 = n11310 & n11311 ;
  assign n11537 = n11533 ^ n11532 ;
  assign n11558 = n11544 ^ n11537 ;
  assign n11308 = n8567 ^ n8503 ;
  assign n11309 = n8568 ^ n8504 ;
  assign n11508 = n11308 & n11309 ;
  assign n11306 = n8565 ^ n8501 ;
  assign n11307 = n8566 ^ n8502 ;
  assign n11507 = n11306 & n11307 ;
  assign n11512 = n11508 ^ n11507 ;
  assign n11304 = n8563 ^ n8499 ;
  assign n11305 = n8564 ^ n8500 ;
  assign n11501 = n11304 & n11305 ;
  assign n11302 = n8561 ^ n8497 ;
  assign n11303 = n8562 ^ n8498 ;
  assign n11500 = n11302 & n11303 ;
  assign n11505 = n11501 ^ n11500 ;
  assign n11526 = n11512 ^ n11505 ;
  assign n11607 = n11558 ^ n11526 ;
  assign n11300 = n8559 ^ n8495 ;
  assign n11301 = n8560 ^ n8496 ;
  assign n11421 = n11300 & n11301 ;
  assign n11298 = n8557 ^ n8493 ;
  assign n11299 = n8558 ^ n8494 ;
  assign n11420 = n11298 & n11299 ;
  assign n11425 = n11421 ^ n11420 ;
  assign n11296 = n8555 ^ n8491 ;
  assign n11297 = n8556 ^ n8492 ;
  assign n11414 = n11296 & n11297 ;
  assign n11294 = n8553 ^ n8489 ;
  assign n11295 = n8554 ^ n8490 ;
  assign n11413 = n11294 & n11295 ;
  assign n11418 = n11414 ^ n11413 ;
  assign n11439 = n11425 ^ n11418 ;
  assign n11292 = n8551 ^ n8487 ;
  assign n11293 = n8552 ^ n8488 ;
  assign n11389 = n11292 & n11293 ;
  assign n11290 = n8549 ^ n8485 ;
  assign n11291 = n8550 ^ n8486 ;
  assign n11388 = n11290 & n11291 ;
  assign n11393 = n11389 ^ n11388 ;
  assign n11288 = n8547 ^ n8483 ;
  assign n11289 = n8548 ^ n8484 ;
  assign n11382 = n11288 & n11289 ;
  assign n11286 = n8545 ^ n8481 ;
  assign n11287 = n8546 ^ n8482 ;
  assign n11381 = n11286 & n11287 ;
  assign n11386 = n11382 ^ n11381 ;
  assign n11407 = n11393 ^ n11386 ;
  assign n11488 = n11439 ^ n11407 ;
  assign n11761 = n11607 ^ n11488 ;
  assign n12640 = n12165 ^ n11761 ;
  assign n12720 = n12688 ^ n12640 ;
  assign n12721 = n12720 ^ n11255 ;
  assign n12912 = n12816 ^ n12721 ;
  assign n8640 = n8450 ^ n8385 ;
  assign n12913 = n12912 ^ n8640 ;
  assign n11945 = n11348 ^ n11346 ;
  assign n11946 = n11349 ^ n11347 ;
  assign n11947 = n11945 & n11946 ;
  assign n11949 = n11947 ^ n11943 ;
  assign n11938 = n11344 ^ n11342 ;
  assign n11939 = n11345 ^ n11343 ;
  assign n11940 = n11938 & n11939 ;
  assign n11942 = n11940 ^ n11936 ;
  assign n11963 = n11949 ^ n11942 ;
  assign n11913 = n11340 ^ n11338 ;
  assign n11914 = n11341 ^ n11339 ;
  assign n11915 = n11913 & n11914 ;
  assign n11917 = n11915 ^ n11911 ;
  assign n11906 = n11336 ^ n11334 ;
  assign n11907 = n11337 ^ n11335 ;
  assign n11908 = n11906 & n11907 ;
  assign n11910 = n11908 ^ n11904 ;
  assign n11931 = n11917 ^ n11910 ;
  assign n12012 = n11963 ^ n11931 ;
  assign n11826 = n11332 ^ n11330 ;
  assign n11827 = n11333 ^ n11331 ;
  assign n11828 = n11826 & n11827 ;
  assign n11830 = n11828 ^ n11824 ;
  assign n11819 = n11328 ^ n11326 ;
  assign n11820 = n11329 ^ n11327 ;
  assign n11821 = n11819 & n11820 ;
  assign n11823 = n11821 ^ n11817 ;
  assign n11844 = n11830 ^ n11823 ;
  assign n11794 = n11324 ^ n11322 ;
  assign n11795 = n11325 ^ n11323 ;
  assign n11796 = n11794 & n11795 ;
  assign n11798 = n11796 ^ n11792 ;
  assign n11787 = n11320 ^ n11318 ;
  assign n11788 = n11321 ^ n11319 ;
  assign n11789 = n11787 & n11788 ;
  assign n11791 = n11789 ^ n11785 ;
  assign n11812 = n11798 ^ n11791 ;
  assign n11893 = n11844 ^ n11812 ;
  assign n12166 = n12012 ^ n11893 ;
  assign n11541 = n11316 ^ n11314 ;
  assign n11542 = n11317 ^ n11315 ;
  assign n11543 = n11541 & n11542 ;
  assign n11545 = n11543 ^ n11539 ;
  assign n11534 = n11312 ^ n11310 ;
  assign n11535 = n11313 ^ n11311 ;
  assign n11536 = n11534 & n11535 ;
  assign n11538 = n11536 ^ n11532 ;
  assign n11559 = n11545 ^ n11538 ;
  assign n11509 = n11308 ^ n11306 ;
  assign n11510 = n11309 ^ n11307 ;
  assign n11511 = n11509 & n11510 ;
  assign n11513 = n11511 ^ n11507 ;
  assign n11502 = n11304 ^ n11302 ;
  assign n11503 = n11305 ^ n11303 ;
  assign n11504 = n11502 & n11503 ;
  assign n11506 = n11504 ^ n11500 ;
  assign n11527 = n11513 ^ n11506 ;
  assign n11608 = n11559 ^ n11527 ;
  assign n11422 = n11300 ^ n11298 ;
  assign n11423 = n11301 ^ n11299 ;
  assign n11424 = n11422 & n11423 ;
  assign n11426 = n11424 ^ n11420 ;
  assign n11415 = n11296 ^ n11294 ;
  assign n11416 = n11297 ^ n11295 ;
  assign n11417 = n11415 & n11416 ;
  assign n11419 = n11417 ^ n11413 ;
  assign n11440 = n11426 ^ n11419 ;
  assign n11390 = n11292 ^ n11290 ;
  assign n11391 = n11293 ^ n11291 ;
  assign n11392 = n11390 & n11391 ;
  assign n11394 = n11392 ^ n11388 ;
  assign n11383 = n11288 ^ n11286 ;
  assign n11384 = n11289 ^ n11287 ;
  assign n11385 = n11383 & n11384 ;
  assign n11387 = n11385 ^ n11381 ;
  assign n11408 = n11394 ^ n11387 ;
  assign n11489 = n11440 ^ n11408 ;
  assign n11762 = n11608 ^ n11489 ;
  assign n12641 = n12166 ^ n11762 ;
  assign n12722 = n12689 ^ n12641 ;
  assign n12723 = n12722 ^ n11257 ;
  assign n12914 = n12817 ^ n12723 ;
  assign n8641 = n8452 ^ n8386 ;
  assign n12915 = n12914 ^ n8641 ;
  assign n11952 = n11348 ^ n11344 ;
  assign n11953 = n11349 ^ n11345 ;
  assign n11956 = n11952 & n11953 ;
  assign n11950 = n11346 ^ n11342 ;
  assign n11951 = n11347 ^ n11343 ;
  assign n11955 = n11950 & n11951 ;
  assign n11960 = n11956 ^ n11955 ;
  assign n11964 = n11962 ^ n11960 ;
  assign n11965 = n11964 ^ n11949 ;
  assign n11920 = n11340 ^ n11336 ;
  assign n11921 = n11341 ^ n11337 ;
  assign n11924 = n11920 & n11921 ;
  assign n11918 = n11338 ^ n11334 ;
  assign n11919 = n11339 ^ n11335 ;
  assign n11923 = n11918 & n11919 ;
  assign n11928 = n11924 ^ n11923 ;
  assign n11932 = n11930 ^ n11928 ;
  assign n11933 = n11932 ^ n11917 ;
  assign n12013 = n11965 ^ n11933 ;
  assign n11833 = n11332 ^ n11328 ;
  assign n11834 = n11333 ^ n11329 ;
  assign n11837 = n11833 & n11834 ;
  assign n11831 = n11330 ^ n11326 ;
  assign n11832 = n11331 ^ n11327 ;
  assign n11836 = n11831 & n11832 ;
  assign n11841 = n11837 ^ n11836 ;
  assign n11845 = n11843 ^ n11841 ;
  assign n11846 = n11845 ^ n11830 ;
  assign n11801 = n11324 ^ n11320 ;
  assign n11802 = n11325 ^ n11321 ;
  assign n11805 = n11801 & n11802 ;
  assign n11799 = n11322 ^ n11318 ;
  assign n11800 = n11323 ^ n11319 ;
  assign n11804 = n11799 & n11800 ;
  assign n11809 = n11805 ^ n11804 ;
  assign n11813 = n11811 ^ n11809 ;
  assign n11814 = n11813 ^ n11798 ;
  assign n11894 = n11846 ^ n11814 ;
  assign n12167 = n12013 ^ n11894 ;
  assign n11548 = n11316 ^ n11312 ;
  assign n11549 = n11317 ^ n11313 ;
  assign n11552 = n11548 & n11549 ;
  assign n11546 = n11314 ^ n11310 ;
  assign n11547 = n11315 ^ n11311 ;
  assign n11551 = n11546 & n11547 ;
  assign n11556 = n11552 ^ n11551 ;
  assign n11560 = n11558 ^ n11556 ;
  assign n11561 = n11560 ^ n11545 ;
  assign n11516 = n11308 ^ n11304 ;
  assign n11517 = n11309 ^ n11305 ;
  assign n11520 = n11516 & n11517 ;
  assign n11514 = n11306 ^ n11302 ;
  assign n11515 = n11307 ^ n11303 ;
  assign n11519 = n11514 & n11515 ;
  assign n11524 = n11520 ^ n11519 ;
  assign n11528 = n11526 ^ n11524 ;
  assign n11529 = n11528 ^ n11513 ;
  assign n11609 = n11561 ^ n11529 ;
  assign n11429 = n11300 ^ n11296 ;
  assign n11430 = n11301 ^ n11297 ;
  assign n11433 = n11429 & n11430 ;
  assign n11427 = n11298 ^ n11294 ;
  assign n11428 = n11299 ^ n11295 ;
  assign n11432 = n11427 & n11428 ;
  assign n11437 = n11433 ^ n11432 ;
  assign n11441 = n11439 ^ n11437 ;
  assign n11442 = n11441 ^ n11426 ;
  assign n11397 = n11292 ^ n11288 ;
  assign n11398 = n11293 ^ n11289 ;
  assign n11401 = n11397 & n11398 ;
  assign n11395 = n11290 ^ n11286 ;
  assign n11396 = n11291 ^ n11287 ;
  assign n11400 = n11395 & n11396 ;
  assign n11405 = n11401 ^ n11400 ;
  assign n11409 = n11407 ^ n11405 ;
  assign n11410 = n11409 ^ n11394 ;
  assign n11490 = n11442 ^ n11410 ;
  assign n11763 = n11609 ^ n11490 ;
  assign n12642 = n12167 ^ n11763 ;
  assign n12724 = n12690 ^ n12642 ;
  assign n12725 = n12724 ^ n11259 ;
  assign n12916 = n12818 ^ n12725 ;
  assign n8642 = n8454 ^ n8387 ;
  assign n12917 = n12916 ^ n8642 ;
  assign n11957 = n11952 ^ n11950 ;
  assign n11958 = n11953 ^ n11951 ;
  assign n11959 = n11957 & n11958 ;
  assign n11961 = n11959 ^ n11955 ;
  assign n11966 = n11963 ^ n11961 ;
  assign n11954 = n11949 ^ n11948 ;
  assign n11967 = n11966 ^ n11954 ;
  assign n11925 = n11920 ^ n11918 ;
  assign n11926 = n11921 ^ n11919 ;
  assign n11927 = n11925 & n11926 ;
  assign n11929 = n11927 ^ n11923 ;
  assign n11934 = n11931 ^ n11929 ;
  assign n11922 = n11917 ^ n11916 ;
  assign n11935 = n11934 ^ n11922 ;
  assign n12014 = n11967 ^ n11935 ;
  assign n11838 = n11833 ^ n11831 ;
  assign n11839 = n11834 ^ n11832 ;
  assign n11840 = n11838 & n11839 ;
  assign n11842 = n11840 ^ n11836 ;
  assign n11847 = n11844 ^ n11842 ;
  assign n11835 = n11830 ^ n11829 ;
  assign n11848 = n11847 ^ n11835 ;
  assign n11806 = n11801 ^ n11799 ;
  assign n11807 = n11802 ^ n11800 ;
  assign n11808 = n11806 & n11807 ;
  assign n11810 = n11808 ^ n11804 ;
  assign n11815 = n11812 ^ n11810 ;
  assign n11803 = n11798 ^ n11797 ;
  assign n11816 = n11815 ^ n11803 ;
  assign n11895 = n11848 ^ n11816 ;
  assign n12168 = n12014 ^ n11895 ;
  assign n11553 = n11548 ^ n11546 ;
  assign n11554 = n11549 ^ n11547 ;
  assign n11555 = n11553 & n11554 ;
  assign n11557 = n11555 ^ n11551 ;
  assign n11562 = n11559 ^ n11557 ;
  assign n11550 = n11545 ^ n11544 ;
  assign n11563 = n11562 ^ n11550 ;
  assign n11521 = n11516 ^ n11514 ;
  assign n11522 = n11517 ^ n11515 ;
  assign n11523 = n11521 & n11522 ;
  assign n11525 = n11523 ^ n11519 ;
  assign n11530 = n11527 ^ n11525 ;
  assign n11518 = n11513 ^ n11512 ;
  assign n11531 = n11530 ^ n11518 ;
  assign n11610 = n11563 ^ n11531 ;
  assign n11434 = n11429 ^ n11427 ;
  assign n11435 = n11430 ^ n11428 ;
  assign n11436 = n11434 & n11435 ;
  assign n11438 = n11436 ^ n11432 ;
  assign n11443 = n11440 ^ n11438 ;
  assign n11431 = n11426 ^ n11425 ;
  assign n11444 = n11443 ^ n11431 ;
  assign n11402 = n11397 ^ n11395 ;
  assign n11403 = n11398 ^ n11396 ;
  assign n11404 = n11402 & n11403 ;
  assign n11406 = n11404 ^ n11400 ;
  assign n11411 = n11408 ^ n11406 ;
  assign n11399 = n11394 ^ n11393 ;
  assign n11412 = n11411 ^ n11399 ;
  assign n11491 = n11444 ^ n11412 ;
  assign n11764 = n11610 ^ n11491 ;
  assign n12643 = n12168 ^ n11764 ;
  assign n12726 = n12691 ^ n12643 ;
  assign n12727 = n12726 ^ n11261 ;
  assign n12918 = n12819 ^ n12727 ;
  assign n8643 = n8456 ^ n8388 ;
  assign n12919 = n12918 ^ n8643 ;
  assign n11974 = n11348 ^ n11340 ;
  assign n11975 = n11349 ^ n11341 ;
  assign n11987 = n11974 & n11975 ;
  assign n11972 = n11346 ^ n11338 ;
  assign n11973 = n11347 ^ n11339 ;
  assign n11986 = n11972 & n11973 ;
  assign n11991 = n11987 ^ n11986 ;
  assign n11970 = n11344 ^ n11336 ;
  assign n11971 = n11345 ^ n11337 ;
  assign n11980 = n11970 & n11971 ;
  assign n11968 = n11342 ^ n11334 ;
  assign n11969 = n11343 ^ n11335 ;
  assign n11979 = n11968 & n11969 ;
  assign n11984 = n11980 ^ n11979 ;
  assign n12005 = n11991 ^ n11984 ;
  assign n12015 = n12011 ^ n12005 ;
  assign n12016 = n12015 ^ n11965 ;
  assign n11855 = n11332 ^ n11324 ;
  assign n11856 = n11333 ^ n11325 ;
  assign n11868 = n11855 & n11856 ;
  assign n11853 = n11330 ^ n11322 ;
  assign n11854 = n11331 ^ n11323 ;
  assign n11867 = n11853 & n11854 ;
  assign n11872 = n11868 ^ n11867 ;
  assign n11851 = n11328 ^ n11320 ;
  assign n11852 = n11329 ^ n11321 ;
  assign n11861 = n11851 & n11852 ;
  assign n11849 = n11326 ^ n11318 ;
  assign n11850 = n11327 ^ n11319 ;
  assign n11860 = n11849 & n11850 ;
  assign n11865 = n11861 ^ n11860 ;
  assign n11886 = n11872 ^ n11865 ;
  assign n11896 = n11892 ^ n11886 ;
  assign n11897 = n11896 ^ n11846 ;
  assign n12169 = n12016 ^ n11897 ;
  assign n11570 = n11316 ^ n11308 ;
  assign n11571 = n11317 ^ n11309 ;
  assign n11583 = n11570 & n11571 ;
  assign n11568 = n11314 ^ n11306 ;
  assign n11569 = n11315 ^ n11307 ;
  assign n11582 = n11568 & n11569 ;
  assign n11587 = n11583 ^ n11582 ;
  assign n11566 = n11312 ^ n11304 ;
  assign n11567 = n11313 ^ n11305 ;
  assign n11576 = n11566 & n11567 ;
  assign n11564 = n11310 ^ n11302 ;
  assign n11565 = n11311 ^ n11303 ;
  assign n11575 = n11564 & n11565 ;
  assign n11580 = n11576 ^ n11575 ;
  assign n11601 = n11587 ^ n11580 ;
  assign n11611 = n11607 ^ n11601 ;
  assign n11612 = n11611 ^ n11561 ;
  assign n11451 = n11300 ^ n11292 ;
  assign n11452 = n11301 ^ n11293 ;
  assign n11464 = n11451 & n11452 ;
  assign n11449 = n11298 ^ n11290 ;
  assign n11450 = n11299 ^ n11291 ;
  assign n11463 = n11449 & n11450 ;
  assign n11468 = n11464 ^ n11463 ;
  assign n11447 = n11296 ^ n11288 ;
  assign n11448 = n11297 ^ n11289 ;
  assign n11457 = n11447 & n11448 ;
  assign n11445 = n11294 ^ n11286 ;
  assign n11446 = n11295 ^ n11287 ;
  assign n11456 = n11445 & n11446 ;
  assign n11461 = n11457 ^ n11456 ;
  assign n11482 = n11468 ^ n11461 ;
  assign n11492 = n11488 ^ n11482 ;
  assign n11493 = n11492 ^ n11442 ;
  assign n11765 = n11612 ^ n11493 ;
  assign n12644 = n12169 ^ n11765 ;
  assign n12728 = n12692 ^ n12644 ;
  assign n12729 = n12728 ^ n11263 ;
  assign n12920 = n12820 ^ n12729 ;
  assign n8644 = n8458 ^ n8389 ;
  assign n12921 = n12920 ^ n8644 ;
  assign n11988 = n11974 ^ n11972 ;
  assign n11989 = n11975 ^ n11973 ;
  assign n11990 = n11988 & n11989 ;
  assign n11992 = n11990 ^ n11986 ;
  assign n11981 = n11970 ^ n11968 ;
  assign n11982 = n11971 ^ n11969 ;
  assign n11983 = n11981 & n11982 ;
  assign n11985 = n11983 ^ n11979 ;
  assign n12006 = n11992 ^ n11985 ;
  assign n12017 = n12012 ^ n12006 ;
  assign n12018 = n12017 ^ n11967 ;
  assign n11869 = n11855 ^ n11853 ;
  assign n11870 = n11856 ^ n11854 ;
  assign n11871 = n11869 & n11870 ;
  assign n11873 = n11871 ^ n11867 ;
  assign n11862 = n11851 ^ n11849 ;
  assign n11863 = n11852 ^ n11850 ;
  assign n11864 = n11862 & n11863 ;
  assign n11866 = n11864 ^ n11860 ;
  assign n11887 = n11873 ^ n11866 ;
  assign n11898 = n11893 ^ n11887 ;
  assign n11899 = n11898 ^ n11848 ;
  assign n12170 = n12018 ^ n11899 ;
  assign n11584 = n11570 ^ n11568 ;
  assign n11585 = n11571 ^ n11569 ;
  assign n11586 = n11584 & n11585 ;
  assign n11588 = n11586 ^ n11582 ;
  assign n11577 = n11566 ^ n11564 ;
  assign n11578 = n11567 ^ n11565 ;
  assign n11579 = n11577 & n11578 ;
  assign n11581 = n11579 ^ n11575 ;
  assign n11602 = n11588 ^ n11581 ;
  assign n11613 = n11608 ^ n11602 ;
  assign n11614 = n11613 ^ n11563 ;
  assign n11465 = n11451 ^ n11449 ;
  assign n11466 = n11452 ^ n11450 ;
  assign n11467 = n11465 & n11466 ;
  assign n11469 = n11467 ^ n11463 ;
  assign n11458 = n11447 ^ n11445 ;
  assign n11459 = n11448 ^ n11446 ;
  assign n11460 = n11458 & n11459 ;
  assign n11462 = n11460 ^ n11456 ;
  assign n11483 = n11469 ^ n11462 ;
  assign n11494 = n11489 ^ n11483 ;
  assign n11495 = n11494 ^ n11444 ;
  assign n11766 = n11614 ^ n11495 ;
  assign n12645 = n12170 ^ n11766 ;
  assign n12730 = n12693 ^ n12645 ;
  assign n12731 = n12730 ^ n11265 ;
  assign n12922 = n12821 ^ n12731 ;
  assign n8645 = n8460 ^ n8390 ;
  assign n12923 = n12922 ^ n8645 ;
  assign n11995 = n11974 ^ n11970 ;
  assign n11996 = n11975 ^ n11971 ;
  assign n11999 = n11995 & n11996 ;
  assign n11993 = n11972 ^ n11968 ;
  assign n11994 = n11973 ^ n11969 ;
  assign n11998 = n11993 & n11994 ;
  assign n12003 = n11999 ^ n11998 ;
  assign n12007 = n12005 ^ n12003 ;
  assign n12008 = n12007 ^ n11992 ;
  assign n12019 = n12013 ^ n12008 ;
  assign n11977 = n11967 ^ n11962 ;
  assign n12020 = n12019 ^ n11977 ;
  assign n11876 = n11855 ^ n11851 ;
  assign n11877 = n11856 ^ n11852 ;
  assign n11880 = n11876 & n11877 ;
  assign n11874 = n11853 ^ n11849 ;
  assign n11875 = n11854 ^ n11850 ;
  assign n11879 = n11874 & n11875 ;
  assign n11884 = n11880 ^ n11879 ;
  assign n11888 = n11886 ^ n11884 ;
  assign n11889 = n11888 ^ n11873 ;
  assign n11900 = n11894 ^ n11889 ;
  assign n11858 = n11848 ^ n11843 ;
  assign n11901 = n11900 ^ n11858 ;
  assign n12171 = n12020 ^ n11901 ;
  assign n11591 = n11570 ^ n11566 ;
  assign n11592 = n11571 ^ n11567 ;
  assign n11595 = n11591 & n11592 ;
  assign n11589 = n11568 ^ n11564 ;
  assign n11590 = n11569 ^ n11565 ;
  assign n11594 = n11589 & n11590 ;
  assign n11599 = n11595 ^ n11594 ;
  assign n11603 = n11601 ^ n11599 ;
  assign n11604 = n11603 ^ n11588 ;
  assign n11615 = n11609 ^ n11604 ;
  assign n11573 = n11563 ^ n11558 ;
  assign n11616 = n11615 ^ n11573 ;
  assign n11472 = n11451 ^ n11447 ;
  assign n11473 = n11452 ^ n11448 ;
  assign n11476 = n11472 & n11473 ;
  assign n11470 = n11449 ^ n11445 ;
  assign n11471 = n11450 ^ n11446 ;
  assign n11475 = n11470 & n11471 ;
  assign n11480 = n11476 ^ n11475 ;
  assign n11484 = n11482 ^ n11480 ;
  assign n11485 = n11484 ^ n11469 ;
  assign n11496 = n11490 ^ n11485 ;
  assign n11454 = n11444 ^ n11439 ;
  assign n11497 = n11496 ^ n11454 ;
  assign n11767 = n11616 ^ n11497 ;
  assign n12646 = n12171 ^ n11767 ;
  assign n12732 = n12694 ^ n12646 ;
  assign n12733 = n12732 ^ n11267 ;
  assign n12924 = n12822 ^ n12733 ;
  assign n8646 = n8462 ^ n8391 ;
  assign n12925 = n12924 ^ n8646 ;
  assign n12000 = n11995 ^ n11993 ;
  assign n12001 = n11996 ^ n11994 ;
  assign n12002 = n12000 & n12001 ;
  assign n12004 = n12002 ^ n11998 ;
  assign n12009 = n12006 ^ n12004 ;
  assign n11997 = n11992 ^ n11991 ;
  assign n12010 = n12009 ^ n11997 ;
  assign n12021 = n12014 ^ n12010 ;
  assign n11976 = n11967 ^ n11965 ;
  assign n11978 = n11976 ^ n11963 ;
  assign n12022 = n12021 ^ n11978 ;
  assign n11881 = n11876 ^ n11874 ;
  assign n11882 = n11877 ^ n11875 ;
  assign n11883 = n11881 & n11882 ;
  assign n11885 = n11883 ^ n11879 ;
  assign n11890 = n11887 ^ n11885 ;
  assign n11878 = n11873 ^ n11872 ;
  assign n11891 = n11890 ^ n11878 ;
  assign n11902 = n11895 ^ n11891 ;
  assign n11857 = n11848 ^ n11846 ;
  assign n11859 = n11857 ^ n11844 ;
  assign n11903 = n11902 ^ n11859 ;
  assign n12172 = n12022 ^ n11903 ;
  assign n11596 = n11591 ^ n11589 ;
  assign n11597 = n11592 ^ n11590 ;
  assign n11598 = n11596 & n11597 ;
  assign n11600 = n11598 ^ n11594 ;
  assign n11605 = n11602 ^ n11600 ;
  assign n11593 = n11588 ^ n11587 ;
  assign n11606 = n11605 ^ n11593 ;
  assign n11617 = n11610 ^ n11606 ;
  assign n11572 = n11563 ^ n11561 ;
  assign n11574 = n11572 ^ n11559 ;
  assign n11618 = n11617 ^ n11574 ;
  assign n11477 = n11472 ^ n11470 ;
  assign n11478 = n11473 ^ n11471 ;
  assign n11479 = n11477 & n11478 ;
  assign n11481 = n11479 ^ n11475 ;
  assign n11486 = n11483 ^ n11481 ;
  assign n11474 = n11469 ^ n11468 ;
  assign n11487 = n11486 ^ n11474 ;
  assign n11498 = n11491 ^ n11487 ;
  assign n11453 = n11444 ^ n11442 ;
  assign n11455 = n11453 ^ n11440 ;
  assign n11499 = n11498 ^ n11455 ;
  assign n11768 = n11618 ^ n11499 ;
  assign n12647 = n12172 ^ n11768 ;
  assign n12734 = n12695 ^ n12647 ;
  assign n12735 = n12734 ^ n11269 ;
  assign n12926 = n12823 ^ n12735 ;
  assign n8647 = n8464 ^ n8392 ;
  assign n12927 = n12926 ^ n8647 ;
  assign n12037 = n11348 ^ n11332 ;
  assign n12038 = n11349 ^ n11333 ;
  assign n12086 = n12037 & n12038 ;
  assign n12035 = n11346 ^ n11330 ;
  assign n12036 = n11347 ^ n11331 ;
  assign n12085 = n12035 & n12036 ;
  assign n12090 = n12086 ^ n12085 ;
  assign n12033 = n11344 ^ n11328 ;
  assign n12034 = n11345 ^ n11329 ;
  assign n12079 = n12033 & n12034 ;
  assign n12031 = n11342 ^ n11326 ;
  assign n12032 = n11343 ^ n11327 ;
  assign n12078 = n12031 & n12032 ;
  assign n12083 = n12079 ^ n12078 ;
  assign n12104 = n12090 ^ n12083 ;
  assign n12029 = n11340 ^ n11324 ;
  assign n12030 = n11341 ^ n11325 ;
  assign n12054 = n12029 & n12030 ;
  assign n12027 = n11338 ^ n11322 ;
  assign n12028 = n11339 ^ n11323 ;
  assign n12053 = n12027 & n12028 ;
  assign n12058 = n12054 ^ n12053 ;
  assign n12025 = n11336 ^ n11320 ;
  assign n12026 = n11337 ^ n11321 ;
  assign n12047 = n12025 & n12026 ;
  assign n12023 = n11334 ^ n11318 ;
  assign n12024 = n11335 ^ n11319 ;
  assign n12046 = n12023 & n12024 ;
  assign n12051 = n12047 ^ n12046 ;
  assign n12072 = n12058 ^ n12051 ;
  assign n12153 = n12104 ^ n12072 ;
  assign n12173 = n12165 ^ n12153 ;
  assign n12174 = n12173 ^ n12016 ;
  assign n11633 = n11316 ^ n11300 ;
  assign n11634 = n11317 ^ n11301 ;
  assign n11682 = n11633 & n11634 ;
  assign n11631 = n11314 ^ n11298 ;
  assign n11632 = n11315 ^ n11299 ;
  assign n11681 = n11631 & n11632 ;
  assign n11686 = n11682 ^ n11681 ;
  assign n11629 = n11312 ^ n11296 ;
  assign n11630 = n11313 ^ n11297 ;
  assign n11675 = n11629 & n11630 ;
  assign n11627 = n11310 ^ n11294 ;
  assign n11628 = n11311 ^ n11295 ;
  assign n11674 = n11627 & n11628 ;
  assign n11679 = n11675 ^ n11674 ;
  assign n11700 = n11686 ^ n11679 ;
  assign n11625 = n11308 ^ n11292 ;
  assign n11626 = n11309 ^ n11293 ;
  assign n11650 = n11625 & n11626 ;
  assign n11623 = n11306 ^ n11290 ;
  assign n11624 = n11307 ^ n11291 ;
  assign n11649 = n11623 & n11624 ;
  assign n11654 = n11650 ^ n11649 ;
  assign n11621 = n11304 ^ n11288 ;
  assign n11622 = n11305 ^ n11289 ;
  assign n11643 = n11621 & n11622 ;
  assign n11619 = n11302 ^ n11286 ;
  assign n11620 = n11303 ^ n11287 ;
  assign n11642 = n11619 & n11620 ;
  assign n11647 = n11643 ^ n11642 ;
  assign n11668 = n11654 ^ n11647 ;
  assign n11749 = n11700 ^ n11668 ;
  assign n11769 = n11761 ^ n11749 ;
  assign n11770 = n11769 ^ n11612 ;
  assign n12648 = n12174 ^ n11770 ;
  assign n12736 = n12696 ^ n12648 ;
  assign n12737 = n12736 ^ n11271 ;
  assign n12928 = n12824 ^ n12737 ;
  assign n8648 = n8466 ^ n8393 ;
  assign n12929 = n12928 ^ n8648 ;
  assign n12087 = n12037 ^ n12035 ;
  assign n12088 = n12038 ^ n12036 ;
  assign n12089 = n12087 & n12088 ;
  assign n12091 = n12089 ^ n12085 ;
  assign n12080 = n12033 ^ n12031 ;
  assign n12081 = n12034 ^ n12032 ;
  assign n12082 = n12080 & n12081 ;
  assign n12084 = n12082 ^ n12078 ;
  assign n12105 = n12091 ^ n12084 ;
  assign n12055 = n12029 ^ n12027 ;
  assign n12056 = n12030 ^ n12028 ;
  assign n12057 = n12055 & n12056 ;
  assign n12059 = n12057 ^ n12053 ;
  assign n12048 = n12025 ^ n12023 ;
  assign n12049 = n12026 ^ n12024 ;
  assign n12050 = n12048 & n12049 ;
  assign n12052 = n12050 ^ n12046 ;
  assign n12073 = n12059 ^ n12052 ;
  assign n12154 = n12105 ^ n12073 ;
  assign n12175 = n12166 ^ n12154 ;
  assign n12176 = n12175 ^ n12018 ;
  assign n11683 = n11633 ^ n11631 ;
  assign n11684 = n11634 ^ n11632 ;
  assign n11685 = n11683 & n11684 ;
  assign n11687 = n11685 ^ n11681 ;
  assign n11676 = n11629 ^ n11627 ;
  assign n11677 = n11630 ^ n11628 ;
  assign n11678 = n11676 & n11677 ;
  assign n11680 = n11678 ^ n11674 ;
  assign n11701 = n11687 ^ n11680 ;
  assign n11651 = n11625 ^ n11623 ;
  assign n11652 = n11626 ^ n11624 ;
  assign n11653 = n11651 & n11652 ;
  assign n11655 = n11653 ^ n11649 ;
  assign n11644 = n11621 ^ n11619 ;
  assign n11645 = n11622 ^ n11620 ;
  assign n11646 = n11644 & n11645 ;
  assign n11648 = n11646 ^ n11642 ;
  assign n11669 = n11655 ^ n11648 ;
  assign n11750 = n11701 ^ n11669 ;
  assign n11771 = n11762 ^ n11750 ;
  assign n11772 = n11771 ^ n11614 ;
  assign n12649 = n12176 ^ n11772 ;
  assign n12738 = n12697 ^ n12649 ;
  assign n12739 = n12738 ^ n11273 ;
  assign n12930 = n12825 ^ n12739 ;
  assign n8649 = n8468 ^ n8394 ;
  assign n12931 = n12930 ^ n8649 ;
  assign n12094 = n12037 ^ n12033 ;
  assign n12095 = n12038 ^ n12034 ;
  assign n12098 = n12094 & n12095 ;
  assign n12092 = n12035 ^ n12031 ;
  assign n12093 = n12036 ^ n12032 ;
  assign n12097 = n12092 & n12093 ;
  assign n12102 = n12098 ^ n12097 ;
  assign n12106 = n12104 ^ n12102 ;
  assign n12107 = n12106 ^ n12091 ;
  assign n12062 = n12029 ^ n12025 ;
  assign n12063 = n12030 ^ n12026 ;
  assign n12066 = n12062 & n12063 ;
  assign n12060 = n12027 ^ n12023 ;
  assign n12061 = n12028 ^ n12024 ;
  assign n12065 = n12060 & n12061 ;
  assign n12070 = n12066 ^ n12065 ;
  assign n12074 = n12072 ^ n12070 ;
  assign n12075 = n12074 ^ n12059 ;
  assign n12155 = n12107 ^ n12075 ;
  assign n12177 = n12167 ^ n12155 ;
  assign n12178 = n12177 ^ n12020 ;
  assign n11690 = n11633 ^ n11629 ;
  assign n11691 = n11634 ^ n11630 ;
  assign n11694 = n11690 & n11691 ;
  assign n11688 = n11631 ^ n11627 ;
  assign n11689 = n11632 ^ n11628 ;
  assign n11693 = n11688 & n11689 ;
  assign n11698 = n11694 ^ n11693 ;
  assign n11702 = n11700 ^ n11698 ;
  assign n11703 = n11702 ^ n11687 ;
  assign n11658 = n11625 ^ n11621 ;
  assign n11659 = n11626 ^ n11622 ;
  assign n11662 = n11658 & n11659 ;
  assign n11656 = n11623 ^ n11619 ;
  assign n11657 = n11624 ^ n11620 ;
  assign n11661 = n11656 & n11657 ;
  assign n11666 = n11662 ^ n11661 ;
  assign n11670 = n11668 ^ n11666 ;
  assign n11671 = n11670 ^ n11655 ;
  assign n11751 = n11703 ^ n11671 ;
  assign n11773 = n11763 ^ n11751 ;
  assign n11774 = n11773 ^ n11616 ;
  assign n12650 = n12178 ^ n11774 ;
  assign n12740 = n12698 ^ n12650 ;
  assign n12741 = n12740 ^ n11275 ;
  assign n12932 = n12826 ^ n12741 ;
  assign n8650 = n8470 ^ n8395 ;
  assign n12933 = n12932 ^ n8650 ;
  assign n12099 = n12094 ^ n12092 ;
  assign n12100 = n12095 ^ n12093 ;
  assign n12101 = n12099 & n12100 ;
  assign n12103 = n12101 ^ n12097 ;
  assign n12108 = n12105 ^ n12103 ;
  assign n12096 = n12091 ^ n12090 ;
  assign n12109 = n12108 ^ n12096 ;
  assign n12067 = n12062 ^ n12060 ;
  assign n12068 = n12063 ^ n12061 ;
  assign n12069 = n12067 & n12068 ;
  assign n12071 = n12069 ^ n12065 ;
  assign n12076 = n12073 ^ n12071 ;
  assign n12064 = n12059 ^ n12058 ;
  assign n12077 = n12076 ^ n12064 ;
  assign n12156 = n12109 ^ n12077 ;
  assign n12179 = n12168 ^ n12156 ;
  assign n12180 = n12179 ^ n12022 ;
  assign n11695 = n11690 ^ n11688 ;
  assign n11696 = n11691 ^ n11689 ;
  assign n11697 = n11695 & n11696 ;
  assign n11699 = n11697 ^ n11693 ;
  assign n11704 = n11701 ^ n11699 ;
  assign n11692 = n11687 ^ n11686 ;
  assign n11705 = n11704 ^ n11692 ;
  assign n11663 = n11658 ^ n11656 ;
  assign n11664 = n11659 ^ n11657 ;
  assign n11665 = n11663 & n11664 ;
  assign n11667 = n11665 ^ n11661 ;
  assign n11672 = n11669 ^ n11667 ;
  assign n11660 = n11655 ^ n11654 ;
  assign n11673 = n11672 ^ n11660 ;
  assign n11752 = n11705 ^ n11673 ;
  assign n11775 = n11764 ^ n11752 ;
  assign n11776 = n11775 ^ n11618 ;
  assign n12651 = n12180 ^ n11776 ;
  assign n12742 = n12699 ^ n12651 ;
  assign n12743 = n12742 ^ n11277 ;
  assign n12934 = n12827 ^ n12743 ;
  assign n8651 = n8472 ^ n8396 ;
  assign n12935 = n12934 ^ n8651 ;
  assign n12116 = n12037 ^ n12029 ;
  assign n12117 = n12038 ^ n12030 ;
  assign n12129 = n12116 & n12117 ;
  assign n12114 = n12035 ^ n12027 ;
  assign n12115 = n12036 ^ n12028 ;
  assign n12128 = n12114 & n12115 ;
  assign n12133 = n12129 ^ n12128 ;
  assign n12112 = n12033 ^ n12025 ;
  assign n12113 = n12034 ^ n12026 ;
  assign n12122 = n12112 & n12113 ;
  assign n12110 = n12031 ^ n12023 ;
  assign n12111 = n12032 ^ n12024 ;
  assign n12121 = n12110 & n12111 ;
  assign n12126 = n12122 ^ n12121 ;
  assign n12147 = n12133 ^ n12126 ;
  assign n12157 = n12153 ^ n12147 ;
  assign n12158 = n12157 ^ n12107 ;
  assign n12181 = n12169 ^ n12158 ;
  assign n12042 = n12020 ^ n12011 ;
  assign n12182 = n12181 ^ n12042 ;
  assign n11712 = n11633 ^ n11625 ;
  assign n11713 = n11634 ^ n11626 ;
  assign n11725 = n11712 & n11713 ;
  assign n11710 = n11631 ^ n11623 ;
  assign n11711 = n11632 ^ n11624 ;
  assign n11724 = n11710 & n11711 ;
  assign n11729 = n11725 ^ n11724 ;
  assign n11708 = n11629 ^ n11621 ;
  assign n11709 = n11630 ^ n11622 ;
  assign n11718 = n11708 & n11709 ;
  assign n11706 = n11627 ^ n11619 ;
  assign n11707 = n11628 ^ n11620 ;
  assign n11717 = n11706 & n11707 ;
  assign n11722 = n11718 ^ n11717 ;
  assign n11743 = n11729 ^ n11722 ;
  assign n11753 = n11749 ^ n11743 ;
  assign n11754 = n11753 ^ n11703 ;
  assign n11777 = n11765 ^ n11754 ;
  assign n11638 = n11616 ^ n11607 ;
  assign n11778 = n11777 ^ n11638 ;
  assign n12652 = n12182 ^ n11778 ;
  assign n12744 = n12700 ^ n12652 ;
  assign n12745 = n12744 ^ n11279 ;
  assign n12936 = n12828 ^ n12745 ;
  assign n8652 = n8474 ^ n8397 ;
  assign n12937 = n12936 ^ n8652 ;
  assign n12130 = n12116 ^ n12114 ;
  assign n12131 = n12117 ^ n12115 ;
  assign n12132 = n12130 & n12131 ;
  assign n12134 = n12132 ^ n12128 ;
  assign n12123 = n12112 ^ n12110 ;
  assign n12124 = n12113 ^ n12111 ;
  assign n12125 = n12123 & n12124 ;
  assign n12127 = n12125 ^ n12121 ;
  assign n12148 = n12134 ^ n12127 ;
  assign n12159 = n12154 ^ n12148 ;
  assign n12160 = n12159 ^ n12109 ;
  assign n12183 = n12170 ^ n12160 ;
  assign n12043 = n12022 ^ n12012 ;
  assign n12184 = n12183 ^ n12043 ;
  assign n11726 = n11712 ^ n11710 ;
  assign n11727 = n11713 ^ n11711 ;
  assign n11728 = n11726 & n11727 ;
  assign n11730 = n11728 ^ n11724 ;
  assign n11719 = n11708 ^ n11706 ;
  assign n11720 = n11709 ^ n11707 ;
  assign n11721 = n11719 & n11720 ;
  assign n11723 = n11721 ^ n11717 ;
  assign n11744 = n11730 ^ n11723 ;
  assign n11755 = n11750 ^ n11744 ;
  assign n11756 = n11755 ^ n11705 ;
  assign n11779 = n11766 ^ n11756 ;
  assign n11639 = n11618 ^ n11608 ;
  assign n11780 = n11779 ^ n11639 ;
  assign n12653 = n12184 ^ n11780 ;
  assign n12746 = n12701 ^ n12653 ;
  assign n12747 = n12746 ^ n11281 ;
  assign n12938 = n12829 ^ n12747 ;
  assign n8653 = n8476 ^ n8398 ;
  assign n12939 = n12938 ^ n8653 ;
  assign n12137 = n12116 ^ n12112 ;
  assign n12138 = n12117 ^ n12113 ;
  assign n12141 = n12137 & n12138 ;
  assign n12135 = n12114 ^ n12110 ;
  assign n12136 = n12115 ^ n12111 ;
  assign n12140 = n12135 & n12136 ;
  assign n12145 = n12141 ^ n12140 ;
  assign n12149 = n12147 ^ n12145 ;
  assign n12150 = n12149 ^ n12134 ;
  assign n12161 = n12155 ^ n12150 ;
  assign n12119 = n12109 ^ n12104 ;
  assign n12162 = n12161 ^ n12119 ;
  assign n12185 = n12171 ^ n12162 ;
  assign n12040 = n12022 ^ n12016 ;
  assign n12044 = n12040 ^ n12013 ;
  assign n12186 = n12185 ^ n12044 ;
  assign n11733 = n11712 ^ n11708 ;
  assign n11734 = n11713 ^ n11709 ;
  assign n11737 = n11733 & n11734 ;
  assign n11731 = n11710 ^ n11706 ;
  assign n11732 = n11711 ^ n11707 ;
  assign n11736 = n11731 & n11732 ;
  assign n11741 = n11737 ^ n11736 ;
  assign n11745 = n11743 ^ n11741 ;
  assign n11746 = n11745 ^ n11730 ;
  assign n11757 = n11751 ^ n11746 ;
  assign n11715 = n11705 ^ n11700 ;
  assign n11758 = n11757 ^ n11715 ;
  assign n11781 = n11767 ^ n11758 ;
  assign n11636 = n11618 ^ n11612 ;
  assign n11640 = n11636 ^ n11609 ;
  assign n11782 = n11781 ^ n11640 ;
  assign n12654 = n12186 ^ n11782 ;
  assign n12748 = n12702 ^ n12654 ;
  assign n12749 = n12748 ^ n11283 ;
  assign n12940 = n12830 ^ n12749 ;
  assign n8654 = n8478 ^ n8399 ;
  assign n12941 = n12940 ^ n8654 ;
  assign n12142 = n12137 ^ n12135 ;
  assign n12143 = n12138 ^ n12136 ;
  assign n12144 = n12142 & n12143 ;
  assign n12146 = n12144 ^ n12140 ;
  assign n12151 = n12148 ^ n12146 ;
  assign n12139 = n12134 ^ n12133 ;
  assign n12152 = n12151 ^ n12139 ;
  assign n12163 = n12156 ^ n12152 ;
  assign n12118 = n12109 ^ n12107 ;
  assign n12120 = n12118 ^ n12105 ;
  assign n12164 = n12163 ^ n12120 ;
  assign n12187 = n12172 ^ n12164 ;
  assign n12039 = n12022 ^ n12020 ;
  assign n12041 = n12039 ^ n12018 ;
  assign n12045 = n12041 ^ n12014 ;
  assign n12188 = n12187 ^ n12045 ;
  assign n11738 = n11733 ^ n11731 ;
  assign n11739 = n11734 ^ n11732 ;
  assign n11740 = n11738 & n11739 ;
  assign n11742 = n11740 ^ n11736 ;
  assign n11747 = n11744 ^ n11742 ;
  assign n11735 = n11730 ^ n11729 ;
  assign n11748 = n11747 ^ n11735 ;
  assign n11759 = n11752 ^ n11748 ;
  assign n11714 = n11705 ^ n11703 ;
  assign n11716 = n11714 ^ n11701 ;
  assign n11760 = n11759 ^ n11716 ;
  assign n11783 = n11768 ^ n11760 ;
  assign n11635 = n11618 ^ n11616 ;
  assign n11637 = n11635 ^ n11614 ;
  assign n11641 = n11637 ^ n11610 ;
  assign n11784 = n11783 ^ n11641 ;
  assign n12655 = n12188 ^ n11784 ;
  assign n12750 = n12703 ^ n12655 ;
  assign n12751 = n12750 ^ n11285 ;
  assign n12942 = n12831 ^ n12751 ;
  assign n8655 = n8480 ^ n8400 ;
  assign n12943 = n12942 ^ n8655 ;
  assign n12219 = n11348 ^ n11316 ;
  assign n12220 = n11349 ^ n11317 ;
  assign n12395 = n12219 & n12220 ;
  assign n12217 = n11346 ^ n11314 ;
  assign n12218 = n11347 ^ n11315 ;
  assign n12394 = n12217 & n12218 ;
  assign n12399 = n12395 ^ n12394 ;
  assign n12215 = n11344 ^ n11312 ;
  assign n12216 = n11345 ^ n11313 ;
  assign n12388 = n12215 & n12216 ;
  assign n12213 = n11342 ^ n11310 ;
  assign n12214 = n11343 ^ n11311 ;
  assign n12387 = n12213 & n12214 ;
  assign n12392 = n12388 ^ n12387 ;
  assign n12413 = n12399 ^ n12392 ;
  assign n12211 = n11340 ^ n11308 ;
  assign n12212 = n11341 ^ n11309 ;
  assign n12363 = n12211 & n12212 ;
  assign n12209 = n11338 ^ n11306 ;
  assign n12210 = n11339 ^ n11307 ;
  assign n12362 = n12209 & n12210 ;
  assign n12367 = n12363 ^ n12362 ;
  assign n12207 = n11336 ^ n11304 ;
  assign n12208 = n11337 ^ n11305 ;
  assign n12356 = n12207 & n12208 ;
  assign n12205 = n11334 ^ n11302 ;
  assign n12206 = n11335 ^ n11303 ;
  assign n12355 = n12205 & n12206 ;
  assign n12360 = n12356 ^ n12355 ;
  assign n12381 = n12367 ^ n12360 ;
  assign n12462 = n12413 ^ n12381 ;
  assign n12203 = n11332 ^ n11300 ;
  assign n12204 = n11333 ^ n11301 ;
  assign n12276 = n12203 & n12204 ;
  assign n12201 = n11330 ^ n11298 ;
  assign n12202 = n11331 ^ n11299 ;
  assign n12275 = n12201 & n12202 ;
  assign n12280 = n12276 ^ n12275 ;
  assign n12199 = n11328 ^ n11296 ;
  assign n12200 = n11329 ^ n11297 ;
  assign n12269 = n12199 & n12200 ;
  assign n12197 = n11326 ^ n11294 ;
  assign n12198 = n11327 ^ n11295 ;
  assign n12268 = n12197 & n12198 ;
  assign n12273 = n12269 ^ n12268 ;
  assign n12294 = n12280 ^ n12273 ;
  assign n12195 = n11324 ^ n11292 ;
  assign n12196 = n11325 ^ n11293 ;
  assign n12244 = n12195 & n12196 ;
  assign n12193 = n11322 ^ n11290 ;
  assign n12194 = n11323 ^ n11291 ;
  assign n12243 = n12193 & n12194 ;
  assign n12248 = n12244 ^ n12243 ;
  assign n12191 = n11320 ^ n11288 ;
  assign n12192 = n11321 ^ n11289 ;
  assign n12237 = n12191 & n12192 ;
  assign n12189 = n11318 ^ n11286 ;
  assign n12190 = n11319 ^ n11287 ;
  assign n12236 = n12189 & n12190 ;
  assign n12241 = n12237 ^ n12236 ;
  assign n12262 = n12248 ^ n12241 ;
  assign n12343 = n12294 ^ n12262 ;
  assign n12616 = n12462 ^ n12343 ;
  assign n12656 = n12640 ^ n12616 ;
  assign n12657 = n12656 ^ n12174 ;
  assign n12752 = n12704 ^ n12657 ;
  assign n11365 = n11271 ^ n11238 ;
  assign n12753 = n12752 ^ n11365 ;
  assign n12944 = n12832 ^ n12753 ;
  assign n8624 = n8466 ^ n8418 ;
  assign n8656 = n8624 ^ n8401 ;
  assign n12945 = n12944 ^ n8656 ;
  assign n12396 = n12219 ^ n12217 ;
  assign n12397 = n12220 ^ n12218 ;
  assign n12398 = n12396 & n12397 ;
  assign n12400 = n12398 ^ n12394 ;
  assign n12389 = n12215 ^ n12213 ;
  assign n12390 = n12216 ^ n12214 ;
  assign n12391 = n12389 & n12390 ;
  assign n12393 = n12391 ^ n12387 ;
  assign n12414 = n12400 ^ n12393 ;
  assign n12364 = n12211 ^ n12209 ;
  assign n12365 = n12212 ^ n12210 ;
  assign n12366 = n12364 & n12365 ;
  assign n12368 = n12366 ^ n12362 ;
  assign n12357 = n12207 ^ n12205 ;
  assign n12358 = n12208 ^ n12206 ;
  assign n12359 = n12357 & n12358 ;
  assign n12361 = n12359 ^ n12355 ;
  assign n12382 = n12368 ^ n12361 ;
  assign n12463 = n12414 ^ n12382 ;
  assign n12277 = n12203 ^ n12201 ;
  assign n12278 = n12204 ^ n12202 ;
  assign n12279 = n12277 & n12278 ;
  assign n12281 = n12279 ^ n12275 ;
  assign n12270 = n12199 ^ n12197 ;
  assign n12271 = n12200 ^ n12198 ;
  assign n12272 = n12270 & n12271 ;
  assign n12274 = n12272 ^ n12268 ;
  assign n12295 = n12281 ^ n12274 ;
  assign n12245 = n12195 ^ n12193 ;
  assign n12246 = n12196 ^ n12194 ;
  assign n12247 = n12245 & n12246 ;
  assign n12249 = n12247 ^ n12243 ;
  assign n12238 = n12191 ^ n12189 ;
  assign n12239 = n12192 ^ n12190 ;
  assign n12240 = n12238 & n12239 ;
  assign n12242 = n12240 ^ n12236 ;
  assign n12263 = n12249 ^ n12242 ;
  assign n12344 = n12295 ^ n12263 ;
  assign n12617 = n12463 ^ n12344 ;
  assign n12658 = n12641 ^ n12617 ;
  assign n12659 = n12658 ^ n12176 ;
  assign n12754 = n12705 ^ n12659 ;
  assign n11366 = n11273 ^ n11239 ;
  assign n12755 = n12754 ^ n11366 ;
  assign n12946 = n12833 ^ n12755 ;
  assign n8625 = n8468 ^ n8420 ;
  assign n8657 = n8625 ^ n8402 ;
  assign n12947 = n12946 ^ n8657 ;
  assign n12403 = n12219 ^ n12215 ;
  assign n12404 = n12220 ^ n12216 ;
  assign n12407 = n12403 & n12404 ;
  assign n12401 = n12217 ^ n12213 ;
  assign n12402 = n12218 ^ n12214 ;
  assign n12406 = n12401 & n12402 ;
  assign n12411 = n12407 ^ n12406 ;
  assign n12415 = n12413 ^ n12411 ;
  assign n12416 = n12415 ^ n12400 ;
  assign n12371 = n12211 ^ n12207 ;
  assign n12372 = n12212 ^ n12208 ;
  assign n12375 = n12371 & n12372 ;
  assign n12369 = n12209 ^ n12205 ;
  assign n12370 = n12210 ^ n12206 ;
  assign n12374 = n12369 & n12370 ;
  assign n12379 = n12375 ^ n12374 ;
  assign n12383 = n12381 ^ n12379 ;
  assign n12384 = n12383 ^ n12368 ;
  assign n12464 = n12416 ^ n12384 ;
  assign n12284 = n12203 ^ n12199 ;
  assign n12285 = n12204 ^ n12200 ;
  assign n12288 = n12284 & n12285 ;
  assign n12282 = n12201 ^ n12197 ;
  assign n12283 = n12202 ^ n12198 ;
  assign n12287 = n12282 & n12283 ;
  assign n12292 = n12288 ^ n12287 ;
  assign n12296 = n12294 ^ n12292 ;
  assign n12297 = n12296 ^ n12281 ;
  assign n12252 = n12195 ^ n12191 ;
  assign n12253 = n12196 ^ n12192 ;
  assign n12256 = n12252 & n12253 ;
  assign n12250 = n12193 ^ n12189 ;
  assign n12251 = n12194 ^ n12190 ;
  assign n12255 = n12250 & n12251 ;
  assign n12260 = n12256 ^ n12255 ;
  assign n12264 = n12262 ^ n12260 ;
  assign n12265 = n12264 ^ n12249 ;
  assign n12345 = n12297 ^ n12265 ;
  assign n12618 = n12464 ^ n12345 ;
  assign n12660 = n12642 ^ n12618 ;
  assign n12661 = n12660 ^ n12178 ;
  assign n12756 = n12706 ^ n12661 ;
  assign n11367 = n11275 ^ n11240 ;
  assign n12757 = n12756 ^ n11367 ;
  assign n12948 = n12834 ^ n12757 ;
  assign n8626 = n8470 ^ n8422 ;
  assign n8658 = n8626 ^ n8403 ;
  assign n12949 = n12948 ^ n8658 ;
  assign n12408 = n12403 ^ n12401 ;
  assign n12409 = n12404 ^ n12402 ;
  assign n12410 = n12408 & n12409 ;
  assign n12412 = n12410 ^ n12406 ;
  assign n12417 = n12414 ^ n12412 ;
  assign n12405 = n12400 ^ n12399 ;
  assign n12418 = n12417 ^ n12405 ;
  assign n12376 = n12371 ^ n12369 ;
  assign n12377 = n12372 ^ n12370 ;
  assign n12378 = n12376 & n12377 ;
  assign n12380 = n12378 ^ n12374 ;
  assign n12385 = n12382 ^ n12380 ;
  assign n12373 = n12368 ^ n12367 ;
  assign n12386 = n12385 ^ n12373 ;
  assign n12465 = n12418 ^ n12386 ;
  assign n12289 = n12284 ^ n12282 ;
  assign n12290 = n12285 ^ n12283 ;
  assign n12291 = n12289 & n12290 ;
  assign n12293 = n12291 ^ n12287 ;
  assign n12298 = n12295 ^ n12293 ;
  assign n12286 = n12281 ^ n12280 ;
  assign n12299 = n12298 ^ n12286 ;
  assign n12257 = n12252 ^ n12250 ;
  assign n12258 = n12253 ^ n12251 ;
  assign n12259 = n12257 & n12258 ;
  assign n12261 = n12259 ^ n12255 ;
  assign n12266 = n12263 ^ n12261 ;
  assign n12254 = n12249 ^ n12248 ;
  assign n12267 = n12266 ^ n12254 ;
  assign n12346 = n12299 ^ n12267 ;
  assign n12619 = n12465 ^ n12346 ;
  assign n12662 = n12643 ^ n12619 ;
  assign n12663 = n12662 ^ n12180 ;
  assign n12758 = n12707 ^ n12663 ;
  assign n11368 = n11277 ^ n11241 ;
  assign n12759 = n12758 ^ n11368 ;
  assign n12950 = n12835 ^ n12759 ;
  assign n8627 = n8472 ^ n8424 ;
  assign n8659 = n8627 ^ n8404 ;
  assign n12951 = n12950 ^ n8659 ;
  assign n12425 = n12219 ^ n12211 ;
  assign n12426 = n12220 ^ n12212 ;
  assign n12438 = n12425 & n12426 ;
  assign n12423 = n12217 ^ n12209 ;
  assign n12424 = n12218 ^ n12210 ;
  assign n12437 = n12423 & n12424 ;
  assign n12442 = n12438 ^ n12437 ;
  assign n12421 = n12215 ^ n12207 ;
  assign n12422 = n12216 ^ n12208 ;
  assign n12431 = n12421 & n12422 ;
  assign n12419 = n12213 ^ n12205 ;
  assign n12420 = n12214 ^ n12206 ;
  assign n12430 = n12419 & n12420 ;
  assign n12435 = n12431 ^ n12430 ;
  assign n12456 = n12442 ^ n12435 ;
  assign n12466 = n12462 ^ n12456 ;
  assign n12467 = n12466 ^ n12416 ;
  assign n12306 = n12203 ^ n12195 ;
  assign n12307 = n12204 ^ n12196 ;
  assign n12319 = n12306 & n12307 ;
  assign n12304 = n12201 ^ n12193 ;
  assign n12305 = n12202 ^ n12194 ;
  assign n12318 = n12304 & n12305 ;
  assign n12323 = n12319 ^ n12318 ;
  assign n12302 = n12199 ^ n12191 ;
  assign n12303 = n12200 ^ n12192 ;
  assign n12312 = n12302 & n12303 ;
  assign n12300 = n12197 ^ n12189 ;
  assign n12301 = n12198 ^ n12190 ;
  assign n12311 = n12300 & n12301 ;
  assign n12316 = n12312 ^ n12311 ;
  assign n12337 = n12323 ^ n12316 ;
  assign n12347 = n12343 ^ n12337 ;
  assign n12348 = n12347 ^ n12297 ;
  assign n12620 = n12467 ^ n12348 ;
  assign n12664 = n12644 ^ n12620 ;
  assign n12665 = n12664 ^ n12182 ;
  assign n12760 = n12708 ^ n12665 ;
  assign n11369 = n11279 ^ n11242 ;
  assign n12761 = n12760 ^ n11369 ;
  assign n12952 = n12836 ^ n12761 ;
  assign n8628 = n8474 ^ n8426 ;
  assign n8660 = n8628 ^ n8405 ;
  assign n12953 = n12952 ^ n8660 ;
  assign n12439 = n12425 ^ n12423 ;
  assign n12440 = n12426 ^ n12424 ;
  assign n12441 = n12439 & n12440 ;
  assign n12443 = n12441 ^ n12437 ;
  assign n12432 = n12421 ^ n12419 ;
  assign n12433 = n12422 ^ n12420 ;
  assign n12434 = n12432 & n12433 ;
  assign n12436 = n12434 ^ n12430 ;
  assign n12457 = n12443 ^ n12436 ;
  assign n12468 = n12463 ^ n12457 ;
  assign n12469 = n12468 ^ n12418 ;
  assign n12320 = n12306 ^ n12304 ;
  assign n12321 = n12307 ^ n12305 ;
  assign n12322 = n12320 & n12321 ;
  assign n12324 = n12322 ^ n12318 ;
  assign n12313 = n12302 ^ n12300 ;
  assign n12314 = n12303 ^ n12301 ;
  assign n12315 = n12313 & n12314 ;
  assign n12317 = n12315 ^ n12311 ;
  assign n12338 = n12324 ^ n12317 ;
  assign n12349 = n12344 ^ n12338 ;
  assign n12350 = n12349 ^ n12299 ;
  assign n12621 = n12469 ^ n12350 ;
  assign n12666 = n12645 ^ n12621 ;
  assign n12667 = n12666 ^ n12184 ;
  assign n12762 = n12709 ^ n12667 ;
  assign n11370 = n11281 ^ n11243 ;
  assign n12763 = n12762 ^ n11370 ;
  assign n12954 = n12837 ^ n12763 ;
  assign n8629 = n8476 ^ n8428 ;
  assign n8661 = n8629 ^ n8406 ;
  assign n12955 = n12954 ^ n8661 ;
  assign n12446 = n12425 ^ n12421 ;
  assign n12447 = n12426 ^ n12422 ;
  assign n12450 = n12446 & n12447 ;
  assign n12444 = n12423 ^ n12419 ;
  assign n12445 = n12424 ^ n12420 ;
  assign n12449 = n12444 & n12445 ;
  assign n12454 = n12450 ^ n12449 ;
  assign n12458 = n12456 ^ n12454 ;
  assign n12459 = n12458 ^ n12443 ;
  assign n12470 = n12464 ^ n12459 ;
  assign n12428 = n12418 ^ n12413 ;
  assign n12471 = n12470 ^ n12428 ;
  assign n12327 = n12306 ^ n12302 ;
  assign n12328 = n12307 ^ n12303 ;
  assign n12331 = n12327 & n12328 ;
  assign n12325 = n12304 ^ n12300 ;
  assign n12326 = n12305 ^ n12301 ;
  assign n12330 = n12325 & n12326 ;
  assign n12335 = n12331 ^ n12330 ;
  assign n12339 = n12337 ^ n12335 ;
  assign n12340 = n12339 ^ n12324 ;
  assign n12351 = n12345 ^ n12340 ;
  assign n12309 = n12299 ^ n12294 ;
  assign n12352 = n12351 ^ n12309 ;
  assign n12622 = n12471 ^ n12352 ;
  assign n12668 = n12646 ^ n12622 ;
  assign n12669 = n12668 ^ n12186 ;
  assign n12764 = n12710 ^ n12669 ;
  assign n11371 = n11283 ^ n11244 ;
  assign n12765 = n12764 ^ n11371 ;
  assign n12956 = n12838 ^ n12765 ;
  assign n8630 = n8478 ^ n8430 ;
  assign n8662 = n8630 ^ n8407 ;
  assign n12957 = n12956 ^ n8662 ;
  assign n12451 = n12446 ^ n12444 ;
  assign n12452 = n12447 ^ n12445 ;
  assign n12453 = n12451 & n12452 ;
  assign n12455 = n12453 ^ n12449 ;
  assign n12460 = n12457 ^ n12455 ;
  assign n12448 = n12443 ^ n12442 ;
  assign n12461 = n12460 ^ n12448 ;
  assign n12472 = n12465 ^ n12461 ;
  assign n12427 = n12418 ^ n12416 ;
  assign n12429 = n12427 ^ n12414 ;
  assign n12473 = n12472 ^ n12429 ;
  assign n12332 = n12327 ^ n12325 ;
  assign n12333 = n12328 ^ n12326 ;
  assign n12334 = n12332 & n12333 ;
  assign n12336 = n12334 ^ n12330 ;
  assign n12341 = n12338 ^ n12336 ;
  assign n12329 = n12324 ^ n12323 ;
  assign n12342 = n12341 ^ n12329 ;
  assign n12353 = n12346 ^ n12342 ;
  assign n12308 = n12299 ^ n12297 ;
  assign n12310 = n12308 ^ n12295 ;
  assign n12354 = n12353 ^ n12310 ;
  assign n12623 = n12473 ^ n12354 ;
  assign n12670 = n12647 ^ n12623 ;
  assign n12671 = n12670 ^ n12188 ;
  assign n12766 = n12711 ^ n12671 ;
  assign n11372 = n11285 ^ n11245 ;
  assign n12767 = n12766 ^ n11372 ;
  assign n12958 = n12839 ^ n12767 ;
  assign n8631 = n8480 ^ n8432 ;
  assign n8663 = n8631 ^ n8408 ;
  assign n12959 = n12958 ^ n8663 ;
  assign n12488 = n12219 ^ n12203 ;
  assign n12489 = n12220 ^ n12204 ;
  assign n12537 = n12488 & n12489 ;
  assign n12486 = n12217 ^ n12201 ;
  assign n12487 = n12218 ^ n12202 ;
  assign n12536 = n12486 & n12487 ;
  assign n12541 = n12537 ^ n12536 ;
  assign n12484 = n12215 ^ n12199 ;
  assign n12485 = n12216 ^ n12200 ;
  assign n12530 = n12484 & n12485 ;
  assign n12482 = n12213 ^ n12197 ;
  assign n12483 = n12214 ^ n12198 ;
  assign n12529 = n12482 & n12483 ;
  assign n12534 = n12530 ^ n12529 ;
  assign n12555 = n12541 ^ n12534 ;
  assign n12480 = n12211 ^ n12195 ;
  assign n12481 = n12212 ^ n12196 ;
  assign n12505 = n12480 & n12481 ;
  assign n12478 = n12209 ^ n12193 ;
  assign n12479 = n12210 ^ n12194 ;
  assign n12504 = n12478 & n12479 ;
  assign n12509 = n12505 ^ n12504 ;
  assign n12476 = n12207 ^ n12191 ;
  assign n12477 = n12208 ^ n12192 ;
  assign n12498 = n12476 & n12477 ;
  assign n12474 = n12205 ^ n12189 ;
  assign n12475 = n12206 ^ n12190 ;
  assign n12497 = n12474 & n12475 ;
  assign n12502 = n12498 ^ n12497 ;
  assign n12523 = n12509 ^ n12502 ;
  assign n12604 = n12555 ^ n12523 ;
  assign n12624 = n12616 ^ n12604 ;
  assign n12625 = n12624 ^ n12467 ;
  assign n12672 = n12648 ^ n12625 ;
  assign n12228 = n12182 ^ n12165 ;
  assign n12673 = n12672 ^ n12228 ;
  assign n12768 = n12712 ^ n12673 ;
  assign n11357 = n11279 ^ n11255 ;
  assign n11373 = n11357 ^ n11246 ;
  assign n12769 = n12768 ^ n11373 ;
  assign n12960 = n12840 ^ n12769 ;
  assign n8616 = n8474 ^ n8450 ;
  assign n8632 = n8616 ^ n8434 ;
  assign n8664 = n8632 ^ n8409 ;
  assign n12961 = n12960 ^ n8664 ;
  assign n12538 = n12488 ^ n12486 ;
  assign n12539 = n12489 ^ n12487 ;
  assign n12540 = n12538 & n12539 ;
  assign n12542 = n12540 ^ n12536 ;
  assign n12531 = n12484 ^ n12482 ;
  assign n12532 = n12485 ^ n12483 ;
  assign n12533 = n12531 & n12532 ;
  assign n12535 = n12533 ^ n12529 ;
  assign n12556 = n12542 ^ n12535 ;
  assign n12506 = n12480 ^ n12478 ;
  assign n12507 = n12481 ^ n12479 ;
  assign n12508 = n12506 & n12507 ;
  assign n12510 = n12508 ^ n12504 ;
  assign n12499 = n12476 ^ n12474 ;
  assign n12500 = n12477 ^ n12475 ;
  assign n12501 = n12499 & n12500 ;
  assign n12503 = n12501 ^ n12497 ;
  assign n12524 = n12510 ^ n12503 ;
  assign n12605 = n12556 ^ n12524 ;
  assign n12626 = n12617 ^ n12605 ;
  assign n12627 = n12626 ^ n12469 ;
  assign n12674 = n12649 ^ n12627 ;
  assign n12229 = n12184 ^ n12166 ;
  assign n12675 = n12674 ^ n12229 ;
  assign n12770 = n12713 ^ n12675 ;
  assign n11358 = n11281 ^ n11257 ;
  assign n11374 = n11358 ^ n11247 ;
  assign n12771 = n12770 ^ n11374 ;
  assign n12962 = n12841 ^ n12771 ;
  assign n8617 = n8476 ^ n8452 ;
  assign n8633 = n8617 ^ n8436 ;
  assign n8665 = n8633 ^ n8410 ;
  assign n12963 = n12962 ^ n8665 ;
  assign n12545 = n12488 ^ n12484 ;
  assign n12546 = n12489 ^ n12485 ;
  assign n12549 = n12545 & n12546 ;
  assign n12543 = n12486 ^ n12482 ;
  assign n12544 = n12487 ^ n12483 ;
  assign n12548 = n12543 & n12544 ;
  assign n12553 = n12549 ^ n12548 ;
  assign n12557 = n12555 ^ n12553 ;
  assign n12558 = n12557 ^ n12542 ;
  assign n12513 = n12480 ^ n12476 ;
  assign n12514 = n12481 ^ n12477 ;
  assign n12517 = n12513 & n12514 ;
  assign n12511 = n12478 ^ n12474 ;
  assign n12512 = n12479 ^ n12475 ;
  assign n12516 = n12511 & n12512 ;
  assign n12521 = n12517 ^ n12516 ;
  assign n12525 = n12523 ^ n12521 ;
  assign n12526 = n12525 ^ n12510 ;
  assign n12606 = n12558 ^ n12526 ;
  assign n12628 = n12618 ^ n12606 ;
  assign n12629 = n12628 ^ n12471 ;
  assign n12676 = n12650 ^ n12629 ;
  assign n12230 = n12186 ^ n12167 ;
  assign n12677 = n12676 ^ n12230 ;
  assign n12772 = n12714 ^ n12677 ;
  assign n11359 = n11283 ^ n11259 ;
  assign n11375 = n11359 ^ n11248 ;
  assign n12773 = n12772 ^ n11375 ;
  assign n12964 = n12842 ^ n12773 ;
  assign n8618 = n8478 ^ n8454 ;
  assign n8634 = n8618 ^ n8438 ;
  assign n8666 = n8634 ^ n8411 ;
  assign n12965 = n12964 ^ n8666 ;
  assign n12550 = n12545 ^ n12543 ;
  assign n12551 = n12546 ^ n12544 ;
  assign n12552 = n12550 & n12551 ;
  assign n12554 = n12552 ^ n12548 ;
  assign n12559 = n12556 ^ n12554 ;
  assign n12547 = n12542 ^ n12541 ;
  assign n12560 = n12559 ^ n12547 ;
  assign n12518 = n12513 ^ n12511 ;
  assign n12519 = n12514 ^ n12512 ;
  assign n12520 = n12518 & n12519 ;
  assign n12522 = n12520 ^ n12516 ;
  assign n12527 = n12524 ^ n12522 ;
  assign n12515 = n12510 ^ n12509 ;
  assign n12528 = n12527 ^ n12515 ;
  assign n12607 = n12560 ^ n12528 ;
  assign n12630 = n12619 ^ n12607 ;
  assign n12631 = n12630 ^ n12473 ;
  assign n12678 = n12651 ^ n12631 ;
  assign n12231 = n12188 ^ n12168 ;
  assign n12679 = n12678 ^ n12231 ;
  assign n12774 = n12715 ^ n12679 ;
  assign n11360 = n11285 ^ n11261 ;
  assign n11376 = n11360 ^ n11249 ;
  assign n12775 = n12774 ^ n11376 ;
  assign n12966 = n12843 ^ n12775 ;
  assign n8619 = n8480 ^ n8456 ;
  assign n8635 = n8619 ^ n8440 ;
  assign n8667 = n8635 ^ n8412 ;
  assign n12967 = n12966 ^ n8667 ;
  assign n12567 = n12488 ^ n12480 ;
  assign n12568 = n12489 ^ n12481 ;
  assign n12580 = n12567 & n12568 ;
  assign n12565 = n12486 ^ n12478 ;
  assign n12566 = n12487 ^ n12479 ;
  assign n12579 = n12565 & n12566 ;
  assign n12584 = n12580 ^ n12579 ;
  assign n12563 = n12484 ^ n12476 ;
  assign n12564 = n12485 ^ n12477 ;
  assign n12573 = n12563 & n12564 ;
  assign n12561 = n12482 ^ n12474 ;
  assign n12562 = n12483 ^ n12475 ;
  assign n12572 = n12561 & n12562 ;
  assign n12577 = n12573 ^ n12572 ;
  assign n12598 = n12584 ^ n12577 ;
  assign n12608 = n12604 ^ n12598 ;
  assign n12609 = n12608 ^ n12558 ;
  assign n12632 = n12620 ^ n12609 ;
  assign n12493 = n12471 ^ n12462 ;
  assign n12633 = n12632 ^ n12493 ;
  assign n12680 = n12652 ^ n12633 ;
  assign n12224 = n12186 ^ n12174 ;
  assign n12232 = n12224 ^ n12169 ;
  assign n12681 = n12680 ^ n12232 ;
  assign n12776 = n12716 ^ n12681 ;
  assign n11353 = n11283 ^ n11271 ;
  assign n11361 = n11353 ^ n11263 ;
  assign n11377 = n11361 ^ n11250 ;
  assign n12777 = n12776 ^ n11377 ;
  assign n12968 = n12844 ^ n12777 ;
  assign n8612 = n8478 ^ n8466 ;
  assign n8620 = n8612 ^ n8458 ;
  assign n8636 = n8620 ^ n8442 ;
  assign n8668 = n8636 ^ n8413 ;
  assign n12969 = n12968 ^ n8668 ;
  assign n12581 = n12567 ^ n12565 ;
  assign n12582 = n12568 ^ n12566 ;
  assign n12583 = n12581 & n12582 ;
  assign n12585 = n12583 ^ n12579 ;
  assign n12574 = n12563 ^ n12561 ;
  assign n12575 = n12564 ^ n12562 ;
  assign n12576 = n12574 & n12575 ;
  assign n12578 = n12576 ^ n12572 ;
  assign n12599 = n12585 ^ n12578 ;
  assign n12610 = n12605 ^ n12599 ;
  assign n12611 = n12610 ^ n12560 ;
  assign n12634 = n12621 ^ n12611 ;
  assign n12494 = n12473 ^ n12463 ;
  assign n12635 = n12634 ^ n12494 ;
  assign n12682 = n12653 ^ n12635 ;
  assign n12225 = n12188 ^ n12176 ;
  assign n12233 = n12225 ^ n12170 ;
  assign n12683 = n12682 ^ n12233 ;
  assign n12778 = n12717 ^ n12683 ;
  assign n11354 = n11285 ^ n11273 ;
  assign n11362 = n11354 ^ n11265 ;
  assign n11378 = n11362 ^ n11251 ;
  assign n12779 = n12778 ^ n11378 ;
  assign n12970 = n12845 ^ n12779 ;
  assign n8613 = n8480 ^ n8468 ;
  assign n8621 = n8613 ^ n8460 ;
  assign n8637 = n8621 ^ n8444 ;
  assign n8669 = n8637 ^ n8414 ;
  assign n12971 = n12970 ^ n8669 ;
  assign n12588 = n12567 ^ n12563 ;
  assign n12589 = n12568 ^ n12564 ;
  assign n12592 = n12588 & n12589 ;
  assign n12586 = n12565 ^ n12561 ;
  assign n12587 = n12566 ^ n12562 ;
  assign n12591 = n12586 & n12587 ;
  assign n12596 = n12592 ^ n12591 ;
  assign n12600 = n12598 ^ n12596 ;
  assign n12601 = n12600 ^ n12585 ;
  assign n12612 = n12606 ^ n12601 ;
  assign n12570 = n12560 ^ n12555 ;
  assign n12613 = n12612 ^ n12570 ;
  assign n12636 = n12622 ^ n12613 ;
  assign n12491 = n12473 ^ n12467 ;
  assign n12495 = n12491 ^ n12464 ;
  assign n12637 = n12636 ^ n12495 ;
  assign n12684 = n12654 ^ n12637 ;
  assign n12222 = n12188 ^ n12182 ;
  assign n12226 = n12222 ^ n12178 ;
  assign n12234 = n12226 ^ n12171 ;
  assign n12685 = n12684 ^ n12234 ;
  assign n12780 = n12718 ^ n12685 ;
  assign n11351 = n11285 ^ n11279 ;
  assign n11355 = n11351 ^ n11275 ;
  assign n11363 = n11355 ^ n11267 ;
  assign n11379 = n11363 ^ n11252 ;
  assign n12781 = n12780 ^ n11379 ;
  assign n12972 = n12846 ^ n12781 ;
  assign n8610 = n8480 ^ n8474 ;
  assign n8614 = n8610 ^ n8470 ;
  assign n8622 = n8614 ^ n8462 ;
  assign n8638 = n8622 ^ n8446 ;
  assign n8670 = n8638 ^ n8415 ;
  assign n12973 = n12972 ^ n8670 ;
  assign n12593 = n12588 ^ n12586 ;
  assign n12594 = n12589 ^ n12587 ;
  assign n12595 = n12593 & n12594 ;
  assign n12597 = n12595 ^ n12591 ;
  assign n12602 = n12599 ^ n12597 ;
  assign n12590 = n12585 ^ n12584 ;
  assign n12603 = n12602 ^ n12590 ;
  assign n12614 = n12607 ^ n12603 ;
  assign n12569 = n12560 ^ n12558 ;
  assign n12571 = n12569 ^ n12556 ;
  assign n12615 = n12614 ^ n12571 ;
  assign n12638 = n12623 ^ n12615 ;
  assign n12490 = n12473 ^ n12471 ;
  assign n12492 = n12490 ^ n12469 ;
  assign n12496 = n12492 ^ n12465 ;
  assign n12639 = n12638 ^ n12496 ;
  assign n12686 = n12655 ^ n12639 ;
  assign n12221 = n12188 ^ n12186 ;
  assign n12223 = n12221 ^ n12184 ;
  assign n12227 = n12223 ^ n12180 ;
  assign n12235 = n12227 ^ n12172 ;
  assign n12687 = n12686 ^ n12235 ;
  assign n12782 = n12719 ^ n12687 ;
  assign n11350 = n11285 ^ n11283 ;
  assign n11352 = n11350 ^ n11281 ;
  assign n11356 = n11352 ^ n11277 ;
  assign n11364 = n11356 ^ n11269 ;
  assign n11380 = n11364 ^ n11253 ;
  assign n12783 = n12782 ^ n11380 ;
  assign n12974 = n12847 ^ n12783 ;
  assign n8609 = n8480 ^ n8478 ;
  assign n8611 = n8609 ^ n8476 ;
  assign n8615 = n8611 ^ n8472 ;
  assign n8623 = n8615 ^ n8464 ;
  assign n8639 = n8623 ^ n8448 ;
  assign n8671 = n8639 ^ n8416 ;
  assign n12975 = n12974 ^ n8671 ;
  assign y0 = n12784 ;
  assign y1 = n12785 ;
  assign y2 = n12786 ;
  assign y3 = n12787 ;
  assign y4 = n12788 ;
  assign y5 = n12789 ;
  assign y6 = n12790 ;
  assign y7 = n12791 ;
  assign y8 = n12792 ;
  assign y9 = n12793 ;
  assign y10 = n12794 ;
  assign y11 = n12795 ;
  assign y12 = n12796 ;
  assign y13 = n12797 ;
  assign y14 = n12798 ;
  assign y15 = n12799 ;
  assign y16 = n12800 ;
  assign y17 = n12801 ;
  assign y18 = n12802 ;
  assign y19 = n12803 ;
  assign y20 = n12804 ;
  assign y21 = n12805 ;
  assign y22 = n12806 ;
  assign y23 = n12807 ;
  assign y24 = n12808 ;
  assign y25 = n12809 ;
  assign y26 = n12810 ;
  assign y27 = n12811 ;
  assign y28 = n12812 ;
  assign y29 = n12813 ;
  assign y30 = n12814 ;
  assign y31 = n12815 ;
  assign y32 = n12816 ;
  assign y33 = n12817 ;
  assign y34 = n12818 ;
  assign y35 = n12819 ;
  assign y36 = n12820 ;
  assign y37 = n12821 ;
  assign y38 = n12822 ;
  assign y39 = n12823 ;
  assign y40 = n12824 ;
  assign y41 = n12825 ;
  assign y42 = n12826 ;
  assign y43 = n12827 ;
  assign y44 = n12828 ;
  assign y45 = n12829 ;
  assign y46 = n12830 ;
  assign y47 = n12831 ;
  assign y48 = n12832 ;
  assign y49 = n12833 ;
  assign y50 = n12834 ;
  assign y51 = n12835 ;
  assign y52 = n12836 ;
  assign y53 = n12837 ;
  assign y54 = n12838 ;
  assign y55 = n12839 ;
  assign y56 = n12840 ;
  assign y57 = n12841 ;
  assign y58 = n12842 ;
  assign y59 = n12843 ;
  assign y60 = n12844 ;
  assign y61 = n12845 ;
  assign y62 = n12846 ;
  assign y63 = n12847 ;
  assign y64 = n12849 ;
  assign y65 = n12851 ;
  assign y66 = n12853 ;
  assign y67 = n12855 ;
  assign y68 = n12857 ;
  assign y69 = n12859 ;
  assign y70 = n12861 ;
  assign y71 = n12863 ;
  assign y72 = n12865 ;
  assign y73 = n12867 ;
  assign y74 = n12869 ;
  assign y75 = n12871 ;
  assign y76 = n12873 ;
  assign y77 = n12875 ;
  assign y78 = n12877 ;
  assign y79 = n12879 ;
  assign y80 = n12881 ;
  assign y81 = n12883 ;
  assign y82 = n12885 ;
  assign y83 = n12887 ;
  assign y84 = n12889 ;
  assign y85 = n12891 ;
  assign y86 = n12893 ;
  assign y87 = n12895 ;
  assign y88 = n12897 ;
  assign y89 = n12899 ;
  assign y90 = n12901 ;
  assign y91 = n12903 ;
  assign y92 = n12905 ;
  assign y93 = n12907 ;
  assign y94 = n12909 ;
  assign y95 = n12911 ;
  assign y96 = n12913 ;
  assign y97 = n12915 ;
  assign y98 = n12917 ;
  assign y99 = n12919 ;
  assign y100 = n12921 ;
  assign y101 = n12923 ;
  assign y102 = n12925 ;
  assign y103 = n12927 ;
  assign y104 = n12929 ;
  assign y105 = n12931 ;
  assign y106 = n12933 ;
  assign y107 = n12935 ;
  assign y108 = n12937 ;
  assign y109 = n12939 ;
  assign y110 = n12941 ;
  assign y111 = n12943 ;
  assign y112 = n12945 ;
  assign y113 = n12947 ;
  assign y114 = n12949 ;
  assign y115 = n12951 ;
  assign y116 = n12953 ;
  assign y117 = n12955 ;
  assign y118 = n12957 ;
  assign y119 = n12959 ;
  assign y120 = n12961 ;
  assign y121 = n12963 ;
  assign y122 = n12965 ;
  assign y123 = n12967 ;
  assign y124 = n12969 ;
  assign y125 = n12971 ;
  assign y126 = n12973 ;
  assign y127 = n12975 ;
endmodule
