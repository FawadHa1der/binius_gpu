// copyrights Fawad Haider
module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 ;
  assign n57 = x7 & x15 ;
  assign n56 = x6 & x14 ;
  assign n61 = n57 ^ n56 ;
  assign n50 = x5 & x13 ;
  assign n49 = x4 & x12 ;
  assign n54 = n50 ^ n49 ;
  assign n75 = n61 ^ n54 ;
  assign n25 = x3 & x11 ;
  assign n24 = x2 & x10 ;
  assign n29 = n25 ^ n24 ;
  assign n18 = x1 & x9 ;
  assign n17 = x0 & x8 ;
  assign n22 = n18 ^ n17 ;
  assign n43 = n29 ^ n22 ;
  assign n124 = n75 ^ n43 ;
  assign n58 = x7 ^ x6 ;
  assign n59 = x15 ^ x14 ;
  assign n60 = n58 & n59 ;
  assign n62 = n60 ^ n56 ;
  assign n51 = x5 ^ x4 ;
  assign n52 = x13 ^ x12 ;
  assign n53 = n51 & n52 ;
  assign n55 = n53 ^ n49 ;
  assign n76 = n62 ^ n55 ;
  assign n26 = x3 ^ x2 ;
  assign n27 = x11 ^ x10 ;
  assign n28 = n26 & n27 ;
  assign n30 = n28 ^ n24 ;
  assign n19 = x1 ^ x0 ;
  assign n20 = x9 ^ x8 ;
  assign n21 = n19 & n20 ;
  assign n23 = n21 ^ n17 ;
  assign n44 = n30 ^ n23 ;
  assign n125 = n76 ^ n44 ;
  assign n65 = x7 ^ x5 ;
  assign n66 = x15 ^ x13 ;
  assign n69 = n65 & n66 ;
  assign n63 = x6 ^ x4 ;
  assign n64 = x14 ^ x12 ;
  assign n68 = n63 & n64 ;
  assign n73 = n69 ^ n68 ;
  assign n77 = n75 ^ n73 ;
  assign n78 = n77 ^ n62 ;
  assign n33 = x3 ^ x1 ;
  assign n34 = x11 ^ x9 ;
  assign n37 = n33 & n34 ;
  assign n31 = x2 ^ x0 ;
  assign n32 = x10 ^ x8 ;
  assign n36 = n31 & n32 ;
  assign n41 = n37 ^ n36 ;
  assign n45 = n43 ^ n41 ;
  assign n46 = n45 ^ n30 ;
  assign n126 = n78 ^ n46 ;
  assign n70 = n65 ^ n63 ;
  assign n71 = n66 ^ n64 ;
  assign n72 = n70 & n71 ;
  assign n74 = n72 ^ n68 ;
  assign n79 = n76 ^ n74 ;
  assign n67 = n62 ^ n61 ;
  assign n80 = n79 ^ n67 ;
  assign n38 = n33 ^ n31 ;
  assign n39 = n34 ^ n32 ;
  assign n40 = n38 & n39 ;
  assign n42 = n40 ^ n36 ;
  assign n47 = n44 ^ n42 ;
  assign n35 = n30 ^ n29 ;
  assign n48 = n47 ^ n35 ;
  assign n127 = n80 ^ n48 ;
  assign n87 = x7 ^ x3 ;
  assign n88 = x15 ^ x11 ;
  assign n100 = n87 & n88 ;
  assign n85 = x6 ^ x2 ;
  assign n86 = x14 ^ x10 ;
  assign n99 = n85 & n86 ;
  assign n104 = n100 ^ n99 ;
  assign n83 = x5 ^ x1 ;
  assign n84 = x13 ^ x9 ;
  assign n93 = n83 & n84 ;
  assign n81 = x4 ^ x0 ;
  assign n82 = x12 ^ x8 ;
  assign n92 = n81 & n82 ;
  assign n97 = n93 ^ n92 ;
  assign n118 = n104 ^ n97 ;
  assign n128 = n124 ^ n118 ;
  assign n129 = n128 ^ n78 ;
  assign n101 = n87 ^ n85 ;
  assign n102 = n88 ^ n86 ;
  assign n103 = n101 & n102 ;
  assign n105 = n103 ^ n99 ;
  assign n94 = n83 ^ n81 ;
  assign n95 = n84 ^ n82 ;
  assign n96 = n94 & n95 ;
  assign n98 = n96 ^ n92 ;
  assign n119 = n105 ^ n98 ;
  assign n130 = n125 ^ n119 ;
  assign n131 = n130 ^ n80 ;
  assign n108 = n87 ^ n83 ;
  assign n109 = n88 ^ n84 ;
  assign n112 = n108 & n109 ;
  assign n106 = n85 ^ n81 ;
  assign n107 = n86 ^ n82 ;
  assign n111 = n106 & n107 ;
  assign n116 = n112 ^ n111 ;
  assign n120 = n118 ^ n116 ;
  assign n121 = n120 ^ n105 ;
  assign n132 = n126 ^ n121 ;
  assign n90 = n80 ^ n75 ;
  assign n133 = n132 ^ n90 ;
  assign n113 = n108 ^ n106 ;
  assign n114 = n109 ^ n107 ;
  assign n115 = n113 & n114 ;
  assign n117 = n115 ^ n111 ;
  assign n122 = n119 ^ n117 ;
  assign n110 = n105 ^ n104 ;
  assign n123 = n122 ^ n110 ;
  assign n134 = n127 ^ n123 ;
  assign n89 = n80 ^ n78 ;
  assign n91 = n89 ^ n76 ;
  assign n135 = n134 ^ n91 ;
  assign y0 = n124 ;
  assign y1 = n125 ;
  assign y2 = n126 ;
  assign y3 = n127 ;
  assign y4 = n129 ;
  assign y5 = n131 ;
  assign y6 = n133 ;
  assign y7 = n135 ;
endmodule
